magic
tech sky130A
magscale 1 2
timestamp 1651007470
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 218974 700884 218980 700936
rect 219032 700924 219038 700936
rect 306374 700924 306380 700936
rect 219032 700896 306380 700924
rect 219032 700884 219038 700896
rect 306374 700884 306380 700896
rect 306432 700884 306438 700936
rect 264974 700816 264980 700868
rect 265032 700856 265038 700868
rect 413646 700856 413652 700868
rect 265032 700828 413652 700856
rect 265032 700816 265038 700828
rect 413646 700816 413652 700828
rect 413704 700816 413710 700868
rect 154114 700748 154120 700800
rect 154172 700788 154178 700800
rect 320174 700788 320180 700800
rect 154172 700760 320180 700788
rect 154172 700748 154178 700760
rect 320174 700748 320180 700760
rect 320232 700748 320238 700800
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 316034 700720 316040 700732
rect 137888 700692 316040 700720
rect 137888 700680 137894 700692
rect 316034 700680 316040 700692
rect 316092 700680 316098 700732
rect 249794 700612 249800 700664
rect 249852 700652 249858 700664
rect 478506 700652 478512 700664
rect 249852 700624 478512 700652
rect 249852 700612 249858 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 89162 700544 89168 700596
rect 89220 700584 89226 700596
rect 335354 700584 335360 700596
rect 89220 700556 335360 700584
rect 89220 700544 89226 700556
rect 335354 700544 335360 700556
rect 335412 700544 335418 700596
rect 72970 700476 72976 700528
rect 73028 700516 73034 700528
rect 329834 700516 329840 700528
rect 73028 700488 329840 700516
rect 73028 700476 73034 700488
rect 329834 700476 329840 700488
rect 329892 700476 329898 700528
rect 235994 700408 236000 700460
rect 236052 700448 236058 700460
rect 543458 700448 543464 700460
rect 236052 700420 543464 700448
rect 236052 700408 236058 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 349154 700380 349160 700392
rect 24360 700352 349160 700380
rect 24360 700340 24366 700352
rect 349154 700340 349160 700352
rect 349212 700340 349218 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 218054 696940 218060 696992
rect 218112 696980 218118 696992
rect 580166 696980 580172 696992
rect 218112 696952 580172 696980
rect 218112 696940 218118 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 353938 683244 353944 683256
rect 3476 683216 353944 683244
rect 3476 683204 3482 683216
rect 353938 683204 353944 683216
rect 353996 683204 354002 683256
rect 222194 683136 222200 683188
rect 222252 683176 222258 683188
rect 580166 683176 580172 683188
rect 222252 683148 580172 683176
rect 222252 683136 222258 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 282914 677220 282920 677272
rect 282972 677260 282978 677272
rect 292850 677260 292856 677272
rect 282972 677232 292856 677260
rect 282972 677220 282978 677232
rect 292850 677220 292856 677232
rect 292908 677220 292914 677272
rect 278866 677152 278872 677204
rect 278924 677192 278930 677204
rect 347774 677192 347780 677204
rect 278924 677164 347780 677192
rect 278924 677152 278930 677164
rect 347774 677152 347780 677164
rect 347832 677152 347838 677204
rect 269482 677084 269488 677136
rect 269540 677124 269546 677136
rect 364334 677124 364340 677136
rect 269540 677096 364340 677124
rect 269540 677084 269546 677096
rect 364334 677084 364340 677096
rect 364392 677084 364398 677136
rect 201494 677016 201500 677068
rect 201552 677056 201558 677068
rect 302234 677056 302240 677068
rect 201552 677028 302240 677056
rect 201552 677016 201558 677028
rect 302234 677016 302240 677028
rect 302292 677016 302298 677068
rect 255314 676948 255320 677000
rect 255372 676988 255378 677000
rect 429194 676988 429200 677000
rect 255372 676960 429200 676988
rect 255372 676948 255378 676960
rect 429194 676948 429200 676960
rect 429252 676948 429258 677000
rect 241514 676880 241520 676932
rect 241572 676920 241578 676932
rect 494054 676920 494060 676932
rect 241572 676892 494060 676920
rect 241572 676880 241578 676892
rect 494054 676880 494060 676892
rect 494112 676880 494118 676932
rect 227162 676812 227168 676864
rect 227220 676852 227226 676864
rect 558914 676852 558920 676864
rect 227220 676824 558920 676852
rect 227220 676812 227226 676824
rect 558914 676812 558920 676824
rect 558972 676812 558978 676864
rect 266354 675724 266360 675776
rect 266412 675764 266418 675776
rect 288434 675764 288440 675776
rect 266412 675736 288440 675764
rect 266412 675724 266418 675736
rect 288434 675724 288440 675736
rect 288492 675724 288498 675776
rect 274450 675656 274456 675708
rect 274508 675696 274514 675708
rect 331214 675696 331220 675708
rect 274508 675668 331220 675696
rect 274508 675656 274514 675668
rect 331214 675656 331220 675668
rect 331272 675656 331278 675708
rect 260650 675588 260656 675640
rect 260708 675628 260714 675640
rect 397454 675628 397460 675640
rect 260708 675600 397460 675628
rect 260708 675588 260714 675600
rect 397454 675588 397460 675600
rect 397512 675588 397518 675640
rect 246666 675520 246672 675572
rect 246724 675560 246730 675572
rect 462314 675560 462320 675572
rect 246724 675532 462320 675560
rect 246724 675520 246730 675532
rect 462314 675520 462320 675532
rect 462372 675520 462378 675572
rect 232682 675452 232688 675504
rect 232740 675492 232746 675504
rect 527174 675492 527180 675504
rect 232740 675464 527180 675492
rect 232740 675452 232746 675464
rect 527174 675452 527180 675464
rect 527232 675452 527238 675504
rect 194962 675384 194968 675436
rect 195020 675424 195026 675436
rect 557166 675424 557172 675436
rect 195020 675396 557172 675424
rect 195020 675384 195026 675396
rect 557166 675384 557172 675396
rect 557224 675384 557230 675436
rect 180702 675316 180708 675368
rect 180760 675356 180766 675368
rect 556982 675356 556988 675368
rect 180760 675328 556988 675356
rect 180760 675316 180766 675328
rect 556982 675316 556988 675328
rect 557040 675316 557046 675368
rect 166810 675248 166816 675300
rect 166868 675288 166874 675300
rect 555970 675288 555976 675300
rect 166868 675260 555976 675288
rect 166868 675248 166874 675260
rect 555970 675248 555976 675260
rect 556028 675248 556034 675300
rect 157242 675180 157248 675232
rect 157300 675220 157306 675232
rect 555878 675220 555884 675232
rect 157300 675192 555884 675220
rect 157300 675180 157306 675192
rect 555878 675180 555884 675192
rect 555936 675180 555942 675232
rect 148042 675112 148048 675164
rect 148100 675152 148106 675164
rect 555786 675152 555792 675164
rect 148100 675124 555792 675152
rect 148100 675112 148106 675124
rect 555786 675112 555792 675124
rect 555844 675112 555850 675164
rect 133782 675044 133788 675096
rect 133840 675084 133846 675096
rect 554590 675084 554596 675096
rect 133840 675056 554596 675084
rect 133840 675044 133846 675056
rect 554590 675044 554596 675056
rect 554648 675044 554654 675096
rect 119890 674976 119896 675028
rect 119948 675016 119954 675028
rect 554406 675016 554412 675028
rect 119948 674988 554412 675016
rect 119948 674976 119954 674988
rect 554406 674976 554412 674988
rect 554464 674976 554470 675028
rect 91738 674908 91744 674960
rect 91796 674948 91802 674960
rect 580166 674948 580172 674960
rect 91796 674920 580172 674948
rect 91796 674908 91802 674920
rect 580166 674908 580172 674920
rect 580224 674908 580230 674960
rect 4890 674840 4896 674892
rect 4948 674880 4954 674892
rect 513742 674880 513748 674892
rect 4948 674852 513748 674880
rect 4948 674840 4954 674852
rect 513742 674840 513748 674852
rect 513800 674840 513806 674892
rect 284202 674364 284208 674416
rect 284260 674404 284266 674416
rect 299474 674404 299480 674416
rect 284260 674376 299480 674404
rect 284260 674364 284266 674376
rect 299474 674364 299480 674376
rect 299532 674364 299538 674416
rect 234614 674296 234620 674348
rect 234672 674336 234678 674348
rect 297726 674336 297732 674348
rect 234672 674308 297732 674336
rect 234672 674296 234678 674308
rect 297726 674296 297732 674308
rect 297784 674296 297790 674348
rect 169754 674228 169760 674280
rect 169812 674268 169818 674280
rect 311894 674268 311900 674280
rect 169812 674240 311900 674268
rect 169812 674228 169818 674240
rect 311894 674228 311900 674240
rect 311952 674228 311958 674280
rect 104894 674160 104900 674212
rect 104952 674200 104958 674212
rect 325878 674200 325884 674212
rect 104952 674172 325884 674200
rect 104952 674160 104958 674172
rect 325878 674160 325884 674172
rect 325936 674160 325942 674212
rect 40034 674092 40040 674144
rect 40092 674132 40098 674144
rect 340046 674132 340052 674144
rect 40092 674104 340052 674132
rect 40092 674092 40098 674104
rect 340046 674092 340052 674104
rect 340104 674092 340110 674144
rect 204162 674024 204168 674076
rect 204220 674064 204226 674076
rect 557350 674064 557356 674076
rect 204220 674036 557356 674064
rect 204220 674024 204226 674036
rect 557350 674024 557356 674036
rect 557408 674024 557414 674076
rect 13906 673956 13912 674008
rect 13964 673996 13970 674008
rect 368566 673996 368572 674008
rect 13964 673968 368572 673996
rect 13964 673956 13970 673968
rect 368566 673956 368572 673968
rect 368624 673956 368630 674008
rect 8938 673888 8944 673940
rect 8996 673928 9002 673940
rect 372798 673928 372804 673940
rect 8996 673900 372804 673928
rect 8996 673888 9002 673900
rect 372798 673888 372804 673900
rect 372856 673888 372862 673940
rect 11790 673820 11796 673872
rect 11848 673860 11854 673872
rect 386966 673860 386972 673872
rect 11848 673832 386972 673860
rect 11848 673820 11854 673832
rect 386966 673820 386972 673832
rect 387024 673820 387030 673872
rect 6362 673752 6368 673804
rect 6420 673792 6426 673804
rect 400950 673792 400956 673804
rect 6420 673764 400956 673792
rect 6420 673752 6426 673764
rect 400950 673752 400956 673764
rect 401008 673752 401014 673804
rect 6270 673684 6276 673736
rect 6328 673724 6334 673736
rect 415486 673724 415492 673736
rect 6328 673696 415492 673724
rect 6328 673684 6334 673696
rect 415486 673684 415492 673696
rect 415544 673684 415550 673736
rect 6178 673616 6184 673668
rect 6236 673656 6242 673668
rect 429194 673656 429200 673668
rect 6236 673628 429200 673656
rect 6236 673616 6242 673628
rect 429194 673616 429200 673628
rect 429252 673616 429258 673668
rect 5442 673548 5448 673600
rect 5500 673588 5506 673600
rect 443270 673588 443276 673600
rect 5500 673560 443276 673588
rect 5500 673548 5506 673560
rect 443270 673548 443276 673560
rect 443328 673548 443334 673600
rect 3878 673480 3884 673532
rect 3936 673520 3942 673532
rect 457438 673520 457444 673532
rect 3936 673492 457444 673520
rect 3936 673480 3942 673492
rect 457438 673480 457444 673492
rect 457496 673480 457502 673532
rect 198734 672936 198740 672988
rect 198792 672976 198798 672988
rect 377582 672976 377588 672988
rect 198792 672948 377588 672976
rect 198792 672936 198798 672948
rect 377582 672936 377588 672948
rect 377640 672936 377646 672988
rect 175918 672868 175924 672920
rect 175976 672908 175982 672920
rect 392026 672908 392032 672920
rect 175976 672880 392032 672908
rect 175976 672868 175982 672880
rect 392026 672868 392032 672880
rect 392084 672868 392090 672920
rect 395430 672868 395436 672920
rect 395488 672908 395494 672920
rect 452654 672908 452660 672920
rect 395488 672880 452660 672908
rect 395488 672868 395494 672880
rect 452654 672868 452660 672880
rect 452712 672868 452718 672920
rect 105722 672800 105728 672852
rect 105780 672840 105786 672852
rect 405734 672840 405740 672852
rect 105780 672812 405740 672840
rect 105780 672800 105786 672812
rect 405734 672800 405740 672812
rect 405792 672800 405798 672852
rect 115106 672732 115112 672784
rect 115164 672772 115170 672784
rect 139486 672772 139492 672784
rect 115164 672744 139492 672772
rect 115164 672732 115170 672744
rect 139486 672732 139492 672744
rect 139544 672732 139550 672784
rect 152826 672732 152832 672784
rect 152884 672772 152890 672784
rect 555694 672772 555700 672784
rect 152884 672744 555700 672772
rect 152884 672732 152890 672744
rect 555694 672732 555700 672744
rect 555752 672732 555758 672784
rect 10318 672664 10324 672716
rect 10376 672704 10382 672716
rect 419718 672704 419724 672716
rect 10376 672676 419724 672704
rect 10376 672664 10382 672676
rect 419718 672664 419724 672676
rect 419776 672664 419782 672716
rect 419810 672664 419816 672716
rect 419868 672704 419874 672716
rect 480806 672704 480812 672716
rect 419868 672676 480812 672704
rect 419868 672664 419874 672676
rect 480806 672664 480812 672676
rect 480864 672664 480870 672716
rect 138658 672596 138664 672648
rect 138716 672636 138722 672648
rect 555602 672636 555608 672648
rect 138716 672608 555608 672636
rect 138716 672596 138722 672608
rect 555602 672596 555608 672608
rect 555660 672596 555666 672648
rect 13078 672528 13084 672580
rect 13136 672568 13142 672580
rect 433886 672568 433892 672580
rect 13136 672540 433892 672568
rect 13136 672528 13142 672540
rect 433886 672528 433892 672540
rect 433944 672528 433950 672580
rect 54202 672460 54208 672512
rect 54260 672500 54266 672512
rect 117958 672500 117964 672512
rect 54260 672472 117964 672500
rect 54260 672460 54266 672472
rect 117958 672460 117964 672472
rect 118016 672460 118022 672512
rect 124674 672460 124680 672512
rect 124732 672500 124738 672512
rect 555510 672500 555516 672512
rect 124732 672472 555516 672500
rect 124732 672460 124738 672472
rect 555510 672460 555516 672472
rect 555568 672460 555574 672512
rect 4706 672392 4712 672444
rect 4764 672432 4770 672444
rect 448054 672432 448060 672444
rect 4764 672404 448060 672432
rect 4764 672392 4770 672404
rect 448054 672392 448060 672404
rect 448112 672392 448118 672444
rect 448146 672392 448152 672444
rect 448204 672432 448210 672444
rect 509234 672432 509240 672444
rect 448204 672404 509240 672432
rect 448204 672392 448210 672404
rect 509234 672392 509240 672404
rect 509292 672392 509298 672444
rect 5350 672324 5356 672376
rect 5408 672364 5414 672376
rect 462314 672364 462320 672376
rect 5408 672336 462320 672364
rect 5408 672324 5414 672336
rect 462314 672324 462320 672336
rect 462372 672324 462378 672376
rect 96338 672256 96344 672308
rect 96396 672296 96402 672308
rect 554130 672296 554136 672308
rect 96396 672268 554136 672296
rect 96396 672256 96402 672268
rect 554130 672256 554136 672268
rect 554188 672256 554194 672308
rect 5258 672188 5264 672240
rect 5316 672228 5322 672240
rect 476206 672228 476212 672240
rect 5316 672200 476212 672228
rect 5316 672188 5322 672200
rect 476206 672188 476212 672200
rect 476264 672188 476270 672240
rect 5166 672120 5172 672172
rect 5224 672160 5230 672172
rect 490190 672160 490196 672172
rect 5224 672132 490196 672160
rect 5224 672120 5230 672132
rect 490190 672120 490196 672132
rect 490248 672120 490254 672172
rect 5074 672052 5080 672104
rect 5132 672092 5138 672104
rect 504358 672092 504364 672104
rect 5132 672064 504364 672092
rect 5132 672052 5138 672064
rect 504358 672052 504364 672064
rect 504416 672052 504422 672104
rect 3326 671508 3332 671560
rect 3384 671548 3390 671560
rect 175918 671548 175924 671560
rect 3384 671520 175924 671548
rect 3384 671508 3390 671520
rect 175918 671508 175924 671520
rect 175976 671508 175982 671560
rect 199746 671508 199752 671560
rect 199804 671548 199810 671560
rect 557258 671548 557264 671560
rect 199804 671520 557264 671548
rect 199804 671508 199810 671520
rect 557258 671508 557264 671520
rect 557316 671508 557322 671560
rect 3234 671440 3240 671492
rect 3292 671480 3298 671492
rect 363414 671480 363420 671492
rect 3292 671452 363420 671480
rect 3292 671440 3298 671452
rect 363414 671440 363420 671452
rect 363472 671440 363478 671492
rect 3050 671372 3056 671424
rect 3108 671412 3114 671424
rect 198734 671412 198740 671424
rect 3108 671384 198740 671412
rect 3108 671372 3114 671384
rect 198734 671372 198740 671384
rect 198792 671372 198798 671424
rect 213730 671372 213736 671424
rect 213788 671412 213794 671424
rect 579614 671412 579620 671424
rect 213788 671384 579620 671412
rect 213788 671372 213794 671384
rect 579614 671372 579620 671384
rect 579672 671372 579678 671424
rect 13354 671304 13360 671356
rect 13412 671344 13418 671356
rect 382274 671344 382280 671356
rect 13412 671316 382280 671344
rect 13412 671304 13418 671316
rect 382274 671304 382280 671316
rect 382332 671304 382338 671356
rect 397086 671304 397092 671356
rect 397144 671344 397150 671356
rect 580534 671344 580540 671356
rect 397144 671316 580540 671344
rect 397144 671304 397150 671316
rect 580534 671304 580540 671316
rect 580592 671304 580598 671356
rect 185578 671236 185584 671288
rect 185636 671276 185642 671288
rect 556062 671276 556068 671288
rect 185636 671248 556068 671276
rect 185636 671236 185642 671248
rect 556062 671236 556068 671248
rect 556120 671236 556126 671288
rect 176194 671168 176200 671220
rect 176252 671208 176258 671220
rect 557074 671208 557080 671220
rect 176252 671180 557080 671208
rect 176252 671168 176258 671180
rect 557074 671168 557080 671180
rect 557132 671168 557138 671220
rect 171594 671100 171600 671152
rect 171652 671140 171658 671152
rect 556890 671140 556896 671152
rect 171652 671112 556896 671140
rect 171652 671100 171658 671112
rect 556890 671100 556896 671112
rect 556948 671100 556954 671152
rect 13262 671032 13268 671084
rect 13320 671072 13326 671084
rect 410334 671072 410340 671084
rect 13320 671044 410340 671072
rect 13320 671032 13326 671044
rect 410334 671032 410340 671044
rect 410392 671032 410398 671084
rect 13170 670964 13176 671016
rect 13228 671004 13234 671016
rect 424502 671004 424508 671016
rect 13228 670976 424508 671004
rect 13228 670964 13234 670976
rect 424502 670964 424508 670976
rect 424560 670964 424566 671016
rect 129274 670896 129280 670948
rect 129332 670936 129338 670948
rect 554498 670936 554504 670948
rect 129332 670908 554504 670936
rect 129332 670896 129338 670908
rect 554498 670896 554504 670908
rect 554556 670896 554562 670948
rect 3786 670828 3792 670880
rect 3844 670868 3850 670880
rect 466822 670868 466828 670880
rect 3844 670840 466828 670868
rect 3844 670828 3850 670840
rect 466822 670828 466828 670840
rect 466880 670828 466886 670880
rect 72970 670760 72976 670812
rect 73028 670800 73034 670812
rect 554038 670800 554044 670812
rect 73028 670772 554044 670800
rect 73028 670760 73034 670772
rect 554038 670760 554044 670772
rect 554096 670760 554102 670812
rect 3418 670692 3424 670744
rect 3476 670732 3482 670744
rect 494974 670732 494980 670744
rect 3476 670704 494980 670732
rect 3476 670692 3482 670704
rect 494974 670692 494980 670704
rect 495032 670692 495038 670744
rect 3970 670216 3976 670268
rect 4028 670256 4034 670268
rect 395430 670256 395436 670268
rect 4028 670228 395436 670256
rect 4028 670216 4034 670228
rect 395430 670216 395436 670228
rect 395488 670216 395494 670268
rect 209130 670148 209136 670200
rect 209188 670188 209194 670200
rect 555326 670188 555332 670200
rect 209188 670160 555332 670188
rect 209188 670148 209194 670160
rect 555326 670148 555332 670160
rect 555384 670148 555390 670200
rect 3602 670080 3608 670132
rect 3660 670120 3666 670132
rect 419810 670120 419816 670132
rect 3660 670092 419816 670120
rect 3660 670080 3666 670092
rect 419810 670080 419816 670092
rect 419868 670080 419874 670132
rect 190178 670012 190184 670064
rect 190236 670052 190242 670064
rect 553946 670052 553952 670064
rect 190236 670024 553952 670052
rect 190236 670012 190242 670024
rect 553946 670012 553952 670024
rect 554004 670012 554010 670064
rect 4062 669944 4068 669996
rect 4120 669984 4126 669996
rect 105722 669984 105728 669996
rect 4120 669956 105728 669984
rect 4120 669944 4126 669956
rect 105722 669944 105728 669956
rect 105780 669944 105786 669996
rect 117958 669944 117964 669996
rect 118016 669984 118022 669996
rect 580350 669984 580356 669996
rect 118016 669956 580356 669984
rect 118016 669944 118022 669956
rect 580350 669944 580356 669956
rect 580408 669944 580414 669996
rect 143442 669876 143448 669928
rect 143500 669916 143506 669928
rect 554682 669916 554688 669928
rect 143500 669888 554688 669916
rect 143500 669876 143506 669888
rect 554682 669876 554688 669888
rect 554740 669876 554746 669928
rect 110322 669808 110328 669860
rect 110380 669848 110386 669860
rect 554222 669848 554228 669860
rect 110380 669820 554228 669848
rect 110380 669808 110386 669820
rect 554222 669808 554228 669820
rect 554280 669808 554286 669860
rect 105722 669740 105728 669792
rect 105780 669780 105786 669792
rect 554314 669780 554320 669792
rect 105780 669752 554320 669780
rect 105780 669740 105786 669752
rect 554314 669740 554320 669752
rect 554372 669740 554378 669792
rect 86862 669672 86868 669724
rect 86920 669712 86926 669724
rect 580902 669712 580908 669724
rect 86920 669684 580908 669712
rect 86920 669672 86926 669684
rect 580902 669672 580908 669684
rect 580960 669672 580966 669724
rect 58802 669604 58808 669656
rect 58860 669644 58866 669656
rect 555418 669644 555424 669656
rect 58860 669616 555424 669644
rect 58860 669604 58866 669616
rect 555418 669604 555424 669616
rect 555476 669604 555482 669656
rect 82354 669536 82360 669588
rect 82412 669576 82418 669588
rect 580718 669576 580724 669588
rect 82412 669548 580724 669576
rect 82412 669536 82418 669548
rect 580718 669536 580724 669548
rect 580776 669536 580782 669588
rect 77570 669468 77576 669520
rect 77628 669508 77634 669520
rect 580810 669508 580816 669520
rect 77628 669480 580816 669508
rect 77628 669468 77634 669480
rect 580810 669468 580816 669480
rect 580868 669468 580874 669520
rect 63402 669400 63408 669452
rect 63460 669440 63466 669452
rect 580626 669440 580632 669452
rect 63460 669412 580632 669440
rect 63460 669400 63466 669412
rect 580626 669400 580632 669412
rect 580684 669400 580690 669452
rect 49418 669332 49424 669384
rect 49476 669372 49482 669384
rect 580442 669372 580448 669384
rect 49476 669344 580448 669372
rect 49476 669332 49482 669344
rect 580442 669332 580448 669344
rect 580500 669332 580506 669384
rect 3142 658180 3148 658232
rect 3200 658220 3206 658232
rect 6454 658220 6460 658232
rect 3200 658192 6460 658220
rect 3200 658180 3206 658192
rect 6454 658180 6460 658192
rect 6512 658180 6518 658232
rect 557350 644376 557356 644428
rect 557408 644416 557414 644428
rect 579982 644416 579988 644428
rect 557408 644388 579988 644416
rect 557408 644376 557414 644388
rect 579982 644376 579988 644388
rect 580040 644376 580046 644428
rect 3142 633360 3148 633412
rect 3200 633400 3206 633412
rect 13814 633400 13820 633412
rect 3200 633372 13820 633400
rect 3200 633360 3206 633372
rect 13814 633360 13820 633372
rect 13872 633360 13878 633412
rect 555326 632000 555332 632052
rect 555384 632040 555390 632052
rect 579982 632040 579988 632052
rect 555384 632012 579988 632040
rect 555384 632000 555390 632012
rect 579982 632000 579988 632012
rect 580040 632000 580046 632052
rect 557258 618196 557264 618248
rect 557316 618236 557322 618248
rect 579982 618236 579988 618248
rect 557316 618208 579988 618236
rect 557316 618196 557322 618208
rect 579982 618196 579988 618208
rect 580040 618196 580046 618248
rect 3142 606772 3148 606824
rect 3200 606812 3206 606824
rect 8938 606812 8944 606824
rect 3200 606784 8944 606812
rect 3200 606772 3206 606784
rect 8938 606772 8944 606784
rect 8996 606772 9002 606824
rect 553946 591948 553952 592000
rect 554004 591988 554010 592000
rect 579798 591988 579804 592000
rect 554004 591960 579804 591988
rect 554004 591948 554010 591960
rect 579798 591948 579804 591960
rect 579856 591948 579862 592000
rect 3234 580932 3240 580984
rect 3292 580972 3298 580984
rect 13354 580972 13360 580984
rect 3292 580944 13360 580972
rect 3292 580932 3298 580944
rect 13354 580932 13360 580944
rect 13412 580932 13418 580984
rect 557166 578144 557172 578196
rect 557224 578184 557230 578196
rect 579798 578184 579804 578196
rect 557224 578156 579804 578184
rect 557224 578144 557230 578156
rect 579798 578144 579804 578156
rect 579856 578144 579862 578196
rect 556062 564340 556068 564392
rect 556120 564380 556126 564392
rect 579982 564380 579988 564392
rect 556120 564352 579988 564380
rect 556120 564340 556126 564352
rect 579982 564340 579988 564352
rect 580040 564340 580046 564392
rect 3326 554684 3332 554736
rect 3384 554724 3390 554736
rect 11790 554724 11796 554736
rect 3384 554696 11796 554724
rect 3384 554684 3390 554696
rect 11790 554684 11796 554696
rect 11848 554684 11854 554736
rect 557074 538160 557080 538212
rect 557132 538200 557138 538212
rect 579982 538200 579988 538212
rect 557132 538172 579988 538200
rect 557132 538160 557138 538172
rect 579982 538160 579988 538172
rect 580040 538160 580046 538212
rect 556982 525716 556988 525768
rect 557040 525756 557046 525768
rect 579982 525756 579988 525768
rect 557040 525728 579988 525756
rect 557040 525716 557046 525728
rect 579982 525716 579988 525728
rect 580040 525716 580046 525768
rect 556890 511912 556896 511964
rect 556948 511952 556954 511964
rect 579982 511952 579988 511964
rect 556948 511924 579988 511952
rect 556948 511912 556954 511924
rect 579982 511912 579988 511924
rect 580040 511912 580046 511964
rect 3234 502120 3240 502172
rect 3292 502160 3298 502172
rect 6362 502160 6368 502172
rect 3292 502132 6368 502160
rect 3292 502120 3298 502132
rect 6362 502120 6368 502132
rect 6420 502120 6426 502172
rect 3326 476008 3332 476060
rect 3384 476048 3390 476060
rect 13262 476048 13268 476060
rect 3384 476020 13268 476048
rect 3384 476008 3390 476020
rect 13262 476008 13268 476020
rect 13320 476008 13326 476060
rect 555970 471928 555976 471980
rect 556028 471968 556034 471980
rect 579798 471968 579804 471980
rect 556028 471940 579804 471968
rect 556028 471928 556034 471940
rect 579798 471928 579804 471940
rect 579856 471928 579862 471980
rect 3326 463632 3332 463684
rect 3384 463672 3390 463684
rect 10318 463672 10324 463684
rect 3384 463644 10324 463672
rect 3384 463632 3390 463644
rect 10318 463632 10324 463644
rect 10376 463632 10382 463684
rect 555878 458124 555884 458176
rect 555936 458164 555942 458176
rect 579982 458164 579988 458176
rect 555936 458136 579988 458164
rect 555936 458124 555942 458136
rect 579982 458124 579988 458136
rect 580040 458124 580046 458176
rect 3142 449556 3148 449608
rect 3200 449596 3206 449608
rect 6270 449596 6276 449608
rect 3200 449568 6276 449596
rect 3200 449556 3206 449568
rect 6270 449556 6276 449568
rect 6328 449556 6334 449608
rect 555786 431876 555792 431928
rect 555844 431916 555850 431928
rect 579982 431916 579988 431928
rect 555844 431888 579988 431916
rect 555844 431876 555850 431888
rect 579982 431876 579988 431888
rect 580040 431876 580046 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 13170 423620 13176 423632
rect 3384 423592 13176 423620
rect 3384 423580 3390 423592
rect 13170 423580 13176 423592
rect 13228 423580 13234 423632
rect 555694 419432 555700 419484
rect 555752 419472 555758 419484
rect 579982 419472 579988 419484
rect 555752 419444 579988 419472
rect 555752 419432 555758 419444
rect 579982 419432 579988 419444
rect 580040 419432 580046 419484
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 13078 411244 13084 411256
rect 3384 411216 13084 411244
rect 3384 411204 3390 411216
rect 13078 411204 13084 411216
rect 13136 411204 13142 411256
rect 554682 405628 554688 405680
rect 554740 405668 554746 405680
rect 579982 405668 579988 405680
rect 554740 405640 579988 405668
rect 554740 405628 554746 405640
rect 579982 405628 579988 405640
rect 580040 405628 580046 405680
rect 3142 398692 3148 398744
rect 3200 398732 3206 398744
rect 6178 398732 6184 398744
rect 3200 398704 6184 398732
rect 3200 398692 3206 398704
rect 6178 398692 6184 398704
rect 6236 398692 6242 398744
rect 554590 379448 554596 379500
rect 554648 379488 554654 379500
rect 579798 379488 579804 379500
rect 554648 379460 579804 379488
rect 554648 379448 554654 379460
rect 579798 379448 579804 379460
rect 579856 379448 579862 379500
rect 555602 365644 555608 365696
rect 555660 365684 555666 365696
rect 579982 365684 579988 365696
rect 555660 365656 579988 365684
rect 555660 365644 555666 365656
rect 579982 365644 579988 365656
rect 580040 365644 580046 365696
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4706 358476 4712 358488
rect 2832 358448 4712 358476
rect 2832 358436 2838 358448
rect 4706 358436 4712 358448
rect 4764 358436 4770 358488
rect 554498 353200 554504 353252
rect 554556 353240 554562 353252
rect 579982 353240 579988 353252
rect 554556 353212 579988 353240
rect 554556 353200 554562 353212
rect 579982 353200 579988 353212
rect 580040 353200 580046 353252
rect 2774 345856 2780 345908
rect 2832 345896 2838 345908
rect 5442 345896 5448 345908
rect 2832 345868 5448 345896
rect 2832 345856 2838 345868
rect 5442 345856 5448 345868
rect 5500 345856 5506 345908
rect 554406 325592 554412 325644
rect 554464 325632 554470 325644
rect 579982 325632 579988 325644
rect 554464 325604 579988 325632
rect 554464 325592 554470 325604
rect 579982 325592 579988 325604
rect 580040 325592 580046 325644
rect 555510 313216 555516 313268
rect 555568 313256 555574 313268
rect 579982 313256 579988 313268
rect 555568 313228 579988 313256
rect 555568 313216 555574 313228
rect 579982 313216 579988 313228
rect 580040 313216 580046 313268
rect 2774 306212 2780 306264
rect 2832 306252 2838 306264
rect 5350 306252 5356 306264
rect 2832 306224 5356 306252
rect 2832 306212 2838 306224
rect 5350 306212 5356 306224
rect 5408 306212 5414 306264
rect 554314 273164 554320 273216
rect 554372 273204 554378 273216
rect 580074 273204 580080 273216
rect 554372 273176 580080 273204
rect 554372 273164 554378 273176
rect 580074 273164 580080 273176
rect 580132 273164 580138 273216
rect 554222 259360 554228 259412
rect 554280 259400 554286 259412
rect 580074 259400 580080 259412
rect 554280 259372 580080 259400
rect 554280 259360 554286 259372
rect 580074 259360 580080 259372
rect 580132 259360 580138 259412
rect 2774 254328 2780 254380
rect 2832 254368 2838 254380
rect 5258 254368 5264 254380
rect 2832 254340 5264 254368
rect 2832 254328 2838 254340
rect 5258 254328 5264 254340
rect 5316 254328 5322 254380
rect 556798 245556 556804 245608
rect 556856 245596 556862 245608
rect 580074 245596 580080 245608
rect 556856 245568 580080 245596
rect 556856 245556 556862 245568
rect 580074 245556 580080 245568
rect 580132 245556 580138 245608
rect 554130 219376 554136 219428
rect 554188 219416 554194 219428
rect 580166 219416 580172 219428
rect 554188 219388 580172 219416
rect 554188 219376 554194 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 2774 202376 2780 202428
rect 2832 202416 2838 202428
rect 5166 202416 5172 202428
rect 2832 202388 5172 202416
rect 2832 202376 2838 202388
rect 5166 202376 5172 202388
rect 5224 202376 5230 202428
rect 554038 166948 554044 167000
rect 554096 166988 554102 167000
rect 579614 166988 579620 167000
rect 554096 166960 579620 166988
rect 554096 166948 554102 166960
rect 579614 166948 579620 166960
rect 579672 166948 579678 167000
rect 2774 149880 2780 149932
rect 2832 149920 2838 149932
rect 5074 149920 5080 149932
rect 2832 149892 5080 149920
rect 2832 149880 2838 149892
rect 5074 149880 5080 149892
rect 5132 149880 5138 149932
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 11698 137952 11704 137964
rect 3292 137924 11704 137952
rect 3292 137912 3298 137924
rect 11698 137912 11704 137924
rect 11756 137912 11762 137964
rect 555418 126896 555424 126948
rect 555476 126936 555482 126948
rect 579614 126936 579620 126948
rect 555476 126908 579620 126936
rect 555476 126896 555482 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 2774 97860 2780 97912
rect 2832 97900 2838 97912
rect 4982 97900 4988 97912
rect 2832 97872 4988 97900
rect 2832 97860 2838 97872
rect 4982 97860 4988 97872
rect 5040 97860 5046 97912
rect 2774 84872 2780 84924
rect 2832 84912 2838 84924
rect 4890 84912 4896 84924
rect 2832 84884 4896 84912
rect 2832 84872 2838 84884
rect 4890 84872 4896 84884
rect 4948 84872 4954 84924
rect 2774 58624 2780 58676
rect 2832 58664 2838 58676
rect 4798 58664 4804 58676
rect 2832 58636 4804 58664
rect 2832 58624 2838 58636
rect 4798 58624 4804 58636
rect 4856 58624 4862 58676
rect 22278 48220 22284 48272
rect 22336 48260 22342 48272
rect 34974 48260 34980 48272
rect 22336 48232 34980 48260
rect 22336 48220 22342 48232
rect 34974 48220 34980 48232
rect 35032 48220 35038 48272
rect 35986 48220 35992 48272
rect 36044 48260 36050 48272
rect 46934 48260 46940 48272
rect 36044 48232 46940 48260
rect 36044 48220 36050 48232
rect 46934 48220 46940 48232
rect 46992 48220 46998 48272
rect 55306 48220 55312 48272
rect 55364 48260 55370 48272
rect 65518 48260 65524 48272
rect 55364 48232 65524 48260
rect 55364 48220 55370 48232
rect 65518 48220 65524 48232
rect 65576 48220 65582 48272
rect 68278 48220 68284 48272
rect 68336 48260 68342 48272
rect 75454 48260 75460 48272
rect 68336 48232 75460 48260
rect 68336 48220 68342 48232
rect 75454 48220 75460 48232
rect 75512 48220 75518 48272
rect 100938 48220 100944 48272
rect 100996 48260 101002 48272
rect 107286 48260 107292 48272
rect 100996 48232 107292 48260
rect 100996 48220 101002 48232
rect 107286 48220 107292 48232
rect 107344 48220 107350 48272
rect 434346 48220 434352 48272
rect 434404 48260 434410 48272
rect 446398 48260 446404 48272
rect 434404 48232 446404 48260
rect 434404 48220 434410 48232
rect 446398 48220 446404 48232
rect 446456 48220 446462 48272
rect 463602 48220 463608 48272
rect 463660 48260 463666 48272
rect 478046 48260 478052 48272
rect 463660 48232 478052 48260
rect 463660 48220 463666 48232
rect 478046 48220 478052 48232
rect 478104 48220 478110 48272
rect 11054 48152 11060 48204
rect 11112 48192 11118 48204
rect 23934 48192 23940 48204
rect 11112 48164 23940 48192
rect 11112 48152 11118 48164
rect 23934 48152 23940 48164
rect 23992 48152 23998 48204
rect 24946 48152 24952 48204
rect 25004 48192 25010 48204
rect 37274 48192 37280 48204
rect 25004 48164 37280 48192
rect 25004 48152 25010 48164
rect 37274 48152 37280 48164
rect 37332 48152 37338 48204
rect 41506 48152 41512 48204
rect 41564 48192 41570 48204
rect 52454 48192 52460 48204
rect 41564 48164 52460 48192
rect 41564 48152 41570 48164
rect 52454 48152 52460 48164
rect 52512 48152 52518 48204
rect 52546 48152 52552 48204
rect 52604 48192 52610 48204
rect 62206 48192 62212 48204
rect 52604 48164 62212 48192
rect 52604 48152 52610 48164
rect 62206 48152 62212 48164
rect 62264 48152 62270 48204
rect 96614 48152 96620 48204
rect 96672 48192 96678 48204
rect 103974 48192 103980 48204
rect 96672 48164 103980 48192
rect 96672 48152 96678 48164
rect 103974 48152 103980 48164
rect 104032 48152 104038 48204
rect 416682 48152 416688 48204
rect 416740 48192 416746 48204
rect 433334 48192 433340 48204
rect 416740 48164 433340 48192
rect 416740 48152 416746 48164
rect 433334 48152 433340 48164
rect 433392 48152 433398 48204
rect 438578 48152 438584 48204
rect 438636 48192 438642 48204
rect 454678 48192 454684 48204
rect 438636 48164 454684 48192
rect 438636 48152 438642 48164
rect 454678 48152 454684 48164
rect 454736 48152 454742 48204
rect 460566 48152 460572 48204
rect 460624 48192 460630 48204
rect 476758 48192 476764 48204
rect 460624 48164 476764 48192
rect 460624 48152 460630 48164
rect 476758 48152 476764 48164
rect 476816 48152 476822 48204
rect 478138 48152 478144 48204
rect 478196 48192 478202 48204
rect 485038 48192 485044 48204
rect 478196 48164 485044 48192
rect 478196 48152 478202 48164
rect 485038 48152 485044 48164
rect 485096 48152 485102 48204
rect 514202 48152 514208 48204
rect 514260 48192 514266 48204
rect 525058 48192 525064 48204
rect 514260 48164 525064 48192
rect 514260 48152 514266 48164
rect 525058 48152 525064 48164
rect 525116 48152 525122 48204
rect 16574 48084 16580 48136
rect 16632 48124 16638 48136
rect 29454 48124 29460 48136
rect 16632 48096 29460 48124
rect 16632 48084 16638 48096
rect 29454 48084 29460 48096
rect 29512 48084 29518 48136
rect 44358 48084 44364 48136
rect 44416 48124 44422 48136
rect 55766 48124 55772 48136
rect 44416 48096 55772 48124
rect 44416 48084 44422 48096
rect 55766 48084 55772 48096
rect 55824 48084 55830 48136
rect 60826 48084 60832 48136
rect 60884 48124 60890 48136
rect 71038 48124 71044 48136
rect 60884 48096 71044 48124
rect 60884 48084 60890 48096
rect 71038 48084 71044 48096
rect 71096 48084 71102 48136
rect 199930 48084 199936 48136
rect 199988 48124 199994 48136
rect 200114 48124 200120 48136
rect 199988 48096 200120 48124
rect 199988 48084 199994 48096
rect 200114 48084 200120 48096
rect 200172 48084 200178 48136
rect 409874 48084 409880 48136
rect 409932 48124 409938 48136
rect 426434 48124 426440 48136
rect 409932 48096 426440 48124
rect 409932 48084 409938 48096
rect 426434 48084 426440 48096
rect 426492 48084 426498 48136
rect 433242 48084 433248 48136
rect 433300 48124 433306 48136
rect 451274 48124 451280 48136
rect 433300 48096 451280 48124
rect 433300 48084 433306 48096
rect 451274 48084 451280 48096
rect 451332 48084 451338 48136
rect 469122 48084 469128 48136
rect 469180 48124 469186 48136
rect 489914 48124 489920 48136
rect 469180 48096 489920 48124
rect 469180 48084 469186 48096
rect 489914 48084 489920 48096
rect 489972 48084 489978 48136
rect 494514 48084 494520 48136
rect 494572 48124 494578 48136
rect 515398 48124 515404 48136
rect 494572 48096 515404 48124
rect 494572 48084 494578 48096
rect 515398 48084 515404 48096
rect 515456 48084 515462 48136
rect 530762 48084 530768 48136
rect 530820 48124 530826 48136
rect 554038 48124 554044 48136
rect 530820 48096 554044 48124
rect 530820 48084 530826 48096
rect 554038 48084 554044 48096
rect 554096 48084 554102 48136
rect 15194 48016 15200 48068
rect 15252 48056 15258 48068
rect 28350 48056 28356 48068
rect 15252 48028 28356 48056
rect 15252 48016 15258 48028
rect 28350 48016 28356 48028
rect 28408 48016 28414 48068
rect 38746 48016 38752 48068
rect 38804 48056 38810 48068
rect 50246 48056 50252 48068
rect 38804 48028 50252 48056
rect 38804 48016 38810 48028
rect 50246 48016 50252 48028
rect 50304 48016 50310 48068
rect 56686 48016 56692 48068
rect 56744 48056 56750 48068
rect 66622 48056 66628 48068
rect 56744 48028 66628 48056
rect 56744 48016 56750 48028
rect 66622 48016 66628 48028
rect 66680 48016 66686 48068
rect 69106 48016 69112 48068
rect 69164 48056 69170 48068
rect 77662 48056 77668 48068
rect 69164 48028 77668 48056
rect 69164 48016 69170 48028
rect 77662 48016 77668 48028
rect 77720 48016 77726 48068
rect 80238 48016 80244 48068
rect 80296 48056 80302 48068
rect 88518 48056 88524 48068
rect 80296 48028 88524 48056
rect 80296 48016 80302 48028
rect 88518 48016 88524 48028
rect 88576 48016 88582 48068
rect 91094 48016 91100 48068
rect 91152 48056 91158 48068
rect 98454 48056 98460 48068
rect 91152 48028 98460 48056
rect 91152 48016 91158 48028
rect 98454 48016 98460 48028
rect 98512 48016 98518 48068
rect 103514 48016 103520 48068
rect 103572 48056 103578 48068
rect 110414 48056 110420 48068
rect 103572 48028 110420 48056
rect 103572 48016 103578 48028
rect 110414 48016 110420 48028
rect 110472 48016 110478 48068
rect 111978 48016 111984 48068
rect 112036 48056 112042 48068
rect 118142 48056 118148 48068
rect 112036 48028 118148 48056
rect 112036 48016 112042 48028
rect 118142 48016 118148 48028
rect 118200 48016 118206 48068
rect 414106 48016 414112 48068
rect 414164 48056 414170 48068
rect 432138 48056 432144 48068
rect 414164 48028 432144 48056
rect 414164 48016 414170 48028
rect 432138 48016 432144 48028
rect 432196 48016 432202 48068
rect 446306 48016 446312 48068
rect 446364 48056 446370 48068
rect 465258 48056 465264 48068
rect 446364 48028 465264 48056
rect 446364 48016 446370 48028
rect 465258 48016 465264 48028
rect 465316 48016 465322 48068
rect 474642 48016 474648 48068
rect 474700 48056 474706 48068
rect 482278 48056 482284 48068
rect 474700 48028 482284 48056
rect 474700 48016 474706 48028
rect 482278 48016 482284 48028
rect 482336 48016 482342 48068
rect 483014 48056 483020 48068
rect 482388 48028 483020 48056
rect 11146 47948 11152 48000
rect 11204 47988 11210 48000
rect 25038 47988 25044 48000
rect 11204 47960 25044 47988
rect 11204 47948 11210 47960
rect 25038 47948 25044 47960
rect 25096 47948 25102 48000
rect 31938 47948 31944 48000
rect 31996 47988 32002 48000
rect 43622 47988 43628 48000
rect 31996 47960 43628 47988
rect 31996 47948 32002 47960
rect 43622 47948 43628 47960
rect 43680 47948 43686 48000
rect 51166 47948 51172 48000
rect 51224 47988 51230 48000
rect 61102 47988 61108 48000
rect 51224 47960 61108 47988
rect 51224 47948 51230 47960
rect 61102 47948 61108 47960
rect 61160 47948 61166 48000
rect 63678 47948 63684 48000
rect 63736 47988 63742 48000
rect 73246 47988 73252 48000
rect 63736 47960 73252 47988
rect 63736 47948 63742 47960
rect 73246 47948 73252 47960
rect 73304 47948 73310 48000
rect 78766 47948 78772 48000
rect 78824 47988 78830 48000
rect 87414 47988 87420 48000
rect 78824 47960 87420 47988
rect 78824 47948 78830 47960
rect 87414 47948 87420 47960
rect 87472 47948 87478 48000
rect 89806 47948 89812 48000
rect 89864 47988 89870 48000
rect 97350 47988 97356 48000
rect 89864 47960 97356 47988
rect 89864 47948 89870 47960
rect 97350 47948 97356 47960
rect 97408 47948 97414 48000
rect 104894 47948 104900 48000
rect 104952 47988 104958 48000
rect 111794 47988 111800 48000
rect 104952 47960 111800 47988
rect 104952 47948 104958 47960
rect 111794 47948 111800 47960
rect 111852 47948 111858 48000
rect 113174 47948 113180 48000
rect 113232 47988 113238 48000
rect 119246 47988 119252 48000
rect 113232 47960 119252 47988
rect 113232 47948 113238 47960
rect 119246 47948 119252 47960
rect 119304 47948 119310 48000
rect 419994 47948 420000 48000
rect 420052 47988 420058 48000
rect 437474 47988 437480 48000
rect 420052 47960 437480 47988
rect 420052 47948 420058 47960
rect 437474 47948 437480 47960
rect 437532 47948 437538 48000
rect 439682 47948 439688 48000
rect 439740 47988 439746 48000
rect 458174 47988 458180 48000
rect 439740 47960 458180 47988
rect 439740 47948 439746 47960
rect 458174 47948 458180 47960
rect 458232 47948 458238 48000
rect 462682 47948 462688 48000
rect 462740 47988 462746 48000
rect 482388 47988 482416 48028
rect 483014 48016 483020 48028
rect 483072 48016 483078 48068
rect 488626 48016 488632 48068
rect 488684 48056 488690 48068
rect 511994 48056 512000 48068
rect 488684 48028 512000 48056
rect 488684 48016 488690 48028
rect 511994 48016 512000 48028
rect 512052 48016 512058 48068
rect 515306 48016 515312 48068
rect 515364 48056 515370 48068
rect 539778 48056 539784 48068
rect 515364 48028 539784 48056
rect 515364 48016 515370 48028
rect 539778 48016 539784 48028
rect 539836 48016 539842 48068
rect 555418 48056 555424 48068
rect 547846 48028 555424 48056
rect 462740 47960 482416 47988
rect 462740 47948 462746 47960
rect 483198 47948 483204 48000
rect 483256 47988 483262 48000
rect 506658 47988 506664 48000
rect 483256 47960 506664 47988
rect 483256 47948 483262 47960
rect 506658 47948 506664 47960
rect 506716 47948 506722 48000
rect 508682 47948 508688 48000
rect 508740 47988 508746 48000
rect 532694 47988 532700 48000
rect 508740 47960 532700 47988
rect 508740 47948 508746 47960
rect 532694 47948 532700 47960
rect 532752 47948 532758 48000
rect 537202 47948 537208 48000
rect 537260 47988 537266 48000
rect 547846 47988 547874 48028
rect 555418 48016 555424 48028
rect 555476 48016 555482 48068
rect 537260 47960 547874 47988
rect 537260 47948 537266 47960
rect 550450 47948 550456 48000
rect 550508 47988 550514 48000
rect 556890 47988 556896 48000
rect 550508 47960 556896 47988
rect 550508 47948 550514 47960
rect 556890 47948 556896 47960
rect 556948 47948 556954 48000
rect 12434 47880 12440 47932
rect 12492 47920 12498 47932
rect 26326 47920 26332 47932
rect 12492 47892 26332 47920
rect 12492 47880 12498 47892
rect 26326 47880 26332 47892
rect 26384 47880 26390 47932
rect 33226 47880 33232 47932
rect 33284 47920 33290 47932
rect 44726 47920 44732 47932
rect 33284 47892 44732 47920
rect 33284 47880 33290 47892
rect 44726 47880 44732 47892
rect 44784 47880 44790 47932
rect 45646 47880 45652 47932
rect 45704 47920 45710 47932
rect 56870 47920 56876 47932
rect 45704 47892 56876 47920
rect 45704 47880 45710 47892
rect 56870 47880 56876 47892
rect 56928 47880 56934 47932
rect 59538 47880 59544 47932
rect 59596 47920 59602 47932
rect 69014 47920 69020 47932
rect 59596 47892 69020 47920
rect 59596 47880 59602 47892
rect 69014 47880 69020 47892
rect 69072 47880 69078 47932
rect 71866 47880 71872 47932
rect 71924 47920 71930 47932
rect 80974 47920 80980 47932
rect 71924 47892 80980 47920
rect 71924 47880 71930 47892
rect 80974 47880 80980 47892
rect 81032 47880 81038 47932
rect 92474 47880 92480 47932
rect 92532 47920 92538 47932
rect 99558 47920 99564 47932
rect 92532 47892 99564 47920
rect 92532 47880 92538 47892
rect 99558 47880 99564 47892
rect 99616 47880 99622 47932
rect 109126 47880 109132 47932
rect 109184 47920 109190 47932
rect 114830 47920 114836 47932
rect 109184 47892 114836 47920
rect 109184 47880 109190 47892
rect 114830 47880 114836 47892
rect 114888 47880 114894 47932
rect 127066 47880 127072 47932
rect 127124 47920 127130 47932
rect 132586 47920 132592 47932
rect 127124 47892 132592 47920
rect 127124 47880 127130 47892
rect 132586 47880 132592 47892
rect 132644 47880 132650 47932
rect 144914 47880 144920 47932
rect 144972 47920 144978 47932
rect 149054 47920 149060 47932
rect 144972 47892 149060 47920
rect 144972 47880 144978 47892
rect 149054 47880 149060 47892
rect 149112 47880 149118 47932
rect 151814 47880 151820 47932
rect 151872 47920 151878 47932
rect 155310 47920 155316 47932
rect 151872 47892 155316 47920
rect 151872 47880 151878 47892
rect 155310 47880 155316 47892
rect 155368 47880 155374 47932
rect 161566 47880 161572 47932
rect 161624 47920 161630 47932
rect 164234 47920 164240 47932
rect 161624 47892 164240 47920
rect 161624 47880 161630 47892
rect 164234 47880 164240 47892
rect 164292 47880 164298 47932
rect 230382 47880 230388 47932
rect 230440 47920 230446 47932
rect 233234 47920 233240 47932
rect 230440 47892 233240 47920
rect 230440 47880 230446 47892
rect 233234 47880 233240 47892
rect 233292 47880 233298 47932
rect 372890 47880 372896 47932
rect 372948 47920 372954 47932
rect 385678 47920 385684 47932
rect 372948 47892 385684 47920
rect 372948 47880 372954 47892
rect 385678 47880 385684 47892
rect 385736 47880 385742 47932
rect 393314 47880 393320 47932
rect 393372 47920 393378 47932
rect 408494 47920 408500 47932
rect 393372 47892 408500 47920
rect 393372 47880 393378 47892
rect 408494 47880 408500 47892
rect 408552 47880 408558 47932
rect 423306 47880 423312 47932
rect 423364 47920 423370 47932
rect 440418 47920 440424 47932
rect 423364 47892 440424 47920
rect 423364 47880 423370 47892
rect 440418 47880 440424 47892
rect 440476 47880 440482 47932
rect 445202 47880 445208 47932
rect 445260 47920 445266 47932
rect 464338 47920 464344 47932
rect 445260 47892 464344 47920
rect 445260 47880 445266 47892
rect 464338 47880 464344 47892
rect 464396 47880 464402 47932
rect 465994 47880 466000 47932
rect 466052 47920 466058 47932
rect 481266 47920 481272 47932
rect 466052 47892 481272 47920
rect 466052 47880 466058 47892
rect 481266 47880 481272 47892
rect 481324 47880 481330 47932
rect 482554 47880 482560 47932
rect 482612 47920 482618 47932
rect 482612 47892 489914 47920
rect 482612 47880 482618 47892
rect 2774 47812 2780 47864
rect 2832 47852 2838 47864
rect 17310 47852 17316 47864
rect 2832 47824 17316 47852
rect 2832 47812 2838 47824
rect 17310 47812 17316 47824
rect 17368 47812 17374 47864
rect 19610 47812 19616 47864
rect 19668 47852 19674 47864
rect 31754 47852 31760 47864
rect 19668 47824 31760 47852
rect 19668 47812 19674 47824
rect 31754 47812 31760 47824
rect 31812 47812 31818 47864
rect 40126 47812 40132 47864
rect 40184 47852 40190 47864
rect 51350 47852 51356 47864
rect 40184 47824 51356 47852
rect 40184 47812 40190 47824
rect 51350 47812 51356 47824
rect 51408 47812 51414 47864
rect 54018 47812 54024 47864
rect 54076 47852 54082 47864
rect 64414 47852 64420 47864
rect 54076 47824 64420 47852
rect 54076 47812 54082 47824
rect 64414 47812 64420 47824
rect 64472 47812 64478 47864
rect 67818 47812 67824 47864
rect 67876 47852 67882 47864
rect 76558 47852 76564 47864
rect 67876 47824 76564 47852
rect 67876 47812 67882 47824
rect 76558 47812 76564 47824
rect 76616 47812 76622 47864
rect 85758 47812 85764 47864
rect 85816 47852 85822 47864
rect 94038 47852 94044 47864
rect 85816 47824 94044 47852
rect 85816 47812 85822 47824
rect 94038 47812 94044 47824
rect 94096 47812 94102 47864
rect 98086 47812 98092 47864
rect 98144 47852 98150 47864
rect 105078 47852 105084 47864
rect 98144 47824 105084 47852
rect 98144 47812 98150 47824
rect 105078 47812 105084 47824
rect 105136 47812 105142 47864
rect 105538 47812 105544 47864
rect 105596 47852 105602 47864
rect 108206 47852 108212 47864
rect 105596 47824 108212 47852
rect 105596 47812 105602 47824
rect 108206 47812 108212 47824
rect 108264 47812 108270 47864
rect 116026 47812 116032 47864
rect 116084 47852 116090 47864
rect 121546 47852 121552 47864
rect 116084 47824 121552 47852
rect 116084 47812 116090 47824
rect 121546 47812 121552 47824
rect 121604 47812 121610 47864
rect 125594 47812 125600 47864
rect 125652 47852 125658 47864
rect 130286 47852 130292 47864
rect 125652 47824 130292 47852
rect 125652 47812 125658 47824
rect 130286 47812 130292 47824
rect 130344 47812 130350 47864
rect 130470 47812 130476 47864
rect 130528 47852 130534 47864
rect 131390 47852 131396 47864
rect 130528 47824 131396 47852
rect 130528 47812 130534 47824
rect 131390 47812 131396 47824
rect 131448 47812 131454 47864
rect 133874 47812 133880 47864
rect 133932 47852 133938 47864
rect 138014 47852 138020 47864
rect 133932 47824 138020 47852
rect 133932 47812 133938 47824
rect 138014 47812 138020 47824
rect 138072 47812 138078 47864
rect 143810 47812 143816 47864
rect 143868 47852 143874 47864
rect 146662 47852 146668 47864
rect 143868 47824 146668 47852
rect 143868 47812 143874 47824
rect 146662 47812 146668 47824
rect 146720 47812 146726 47864
rect 153378 47812 153384 47864
rect 153436 47852 153442 47864
rect 156414 47852 156420 47864
rect 153436 47824 156420 47852
rect 153436 47812 153442 47824
rect 156414 47812 156420 47824
rect 156472 47812 156478 47864
rect 157426 47812 157432 47864
rect 157484 47852 157490 47864
rect 160186 47852 160192 47864
rect 157484 47824 160192 47852
rect 157484 47812 157490 47824
rect 160186 47812 160192 47824
rect 160244 47812 160250 47864
rect 186314 47812 186320 47864
rect 186372 47852 186378 47864
rect 187142 47852 187148 47864
rect 186372 47824 187148 47852
rect 186372 47812 186378 47824
rect 187142 47812 187148 47824
rect 187200 47812 187206 47864
rect 201586 47812 201592 47864
rect 201644 47852 201650 47864
rect 202414 47852 202420 47864
rect 201644 47824 202420 47852
rect 201644 47812 201650 47824
rect 202414 47812 202420 47824
rect 202472 47812 202478 47864
rect 211890 47812 211896 47864
rect 211948 47852 211954 47864
rect 212534 47852 212540 47864
rect 211948 47824 212540 47852
rect 211948 47812 211954 47824
rect 212534 47812 212540 47824
rect 212592 47812 212598 47864
rect 212994 47812 213000 47864
rect 213052 47852 213058 47864
rect 213914 47852 213920 47864
rect 213052 47824 213920 47852
rect 213052 47812 213058 47824
rect 213914 47812 213920 47824
rect 213972 47812 213978 47864
rect 226058 47812 226064 47864
rect 226116 47852 226122 47864
rect 227714 47852 227720 47864
rect 226116 47824 227720 47852
rect 226116 47812 226122 47824
rect 227714 47812 227720 47824
rect 227772 47812 227778 47864
rect 229370 47812 229376 47864
rect 229428 47852 229434 47864
rect 231854 47852 231860 47864
rect 229428 47824 231860 47852
rect 229428 47812 229434 47824
rect 231854 47812 231860 47824
rect 231912 47812 231918 47864
rect 244274 47812 244280 47864
rect 244332 47852 244338 47864
rect 245286 47852 245292 47864
rect 244332 47824 245292 47852
rect 244332 47812 244338 47824
rect 245286 47812 245292 47824
rect 245344 47812 245350 47864
rect 255314 47812 255320 47864
rect 255372 47852 255378 47864
rect 256142 47852 256148 47864
rect 255372 47824 256148 47852
rect 255372 47812 255378 47824
rect 256142 47812 256148 47824
rect 256200 47812 256206 47864
rect 262122 47812 262128 47864
rect 262180 47852 262186 47864
rect 264238 47852 264244 47864
rect 262180 47824 264244 47852
rect 262180 47812 262186 47824
rect 264238 47812 264244 47824
rect 264296 47812 264302 47864
rect 271874 47812 271880 47864
rect 271932 47852 271938 47864
rect 277394 47852 277400 47864
rect 271932 47824 277400 47852
rect 271932 47812 271938 47824
rect 277394 47812 277400 47824
rect 277452 47812 277458 47864
rect 287054 47812 287060 47864
rect 287112 47852 287118 47864
rect 287974 47852 287980 47864
rect 287112 47824 287980 47852
rect 287112 47812 287118 47824
rect 287974 47812 287980 47824
rect 288032 47812 288038 47864
rect 308030 47812 308036 47864
rect 308088 47852 308094 47864
rect 309778 47852 309784 47864
rect 308088 47824 309784 47852
rect 308088 47812 308094 47824
rect 309778 47812 309784 47824
rect 309836 47812 309842 47864
rect 313274 47812 313280 47864
rect 313332 47852 313338 47864
rect 314286 47852 314292 47864
rect 313332 47824 314292 47852
rect 313332 47812 313338 47824
rect 314286 47812 314292 47824
rect 314344 47812 314350 47864
rect 320082 47812 320088 47864
rect 320140 47852 320146 47864
rect 323578 47852 323584 47864
rect 320140 47824 323584 47852
rect 320140 47812 320146 47824
rect 323578 47812 323584 47824
rect 323636 47812 323642 47864
rect 329834 47812 329840 47864
rect 329892 47852 329898 47864
rect 330662 47852 330668 47864
rect 329892 47824 330668 47852
rect 329892 47812 329898 47824
rect 330662 47812 330668 47824
rect 330720 47812 330726 47864
rect 370682 47812 370688 47864
rect 370740 47852 370746 47864
rect 383654 47852 383660 47864
rect 370740 47824 383660 47852
rect 370740 47812 370746 47824
rect 383654 47812 383660 47824
rect 383712 47812 383718 47864
rect 387242 47812 387248 47864
rect 387300 47852 387306 47864
rect 401594 47852 401600 47864
rect 387300 47824 401600 47852
rect 387300 47812 387306 47824
rect 401594 47812 401600 47824
rect 401652 47812 401658 47864
rect 405642 47812 405648 47864
rect 405700 47852 405706 47864
rect 411898 47852 411904 47864
rect 405700 47824 411904 47852
rect 405700 47812 405706 47824
rect 411898 47812 411904 47824
rect 411956 47812 411962 47864
rect 413554 47812 413560 47864
rect 413612 47852 413618 47864
rect 430574 47852 430580 47864
rect 413612 47824 430580 47852
rect 413612 47812 413618 47824
rect 430574 47812 430580 47824
rect 430632 47812 430638 47864
rect 436554 47812 436560 47864
rect 436612 47852 436618 47864
rect 455414 47852 455420 47864
rect 436612 47824 455420 47852
rect 436612 47812 436618 47824
rect 455414 47812 455420 47824
rect 455472 47812 455478 47864
rect 456886 47812 456892 47864
rect 456944 47852 456950 47864
rect 457806 47852 457812 47864
rect 456944 47824 457812 47852
rect 456944 47812 456950 47824
rect 457806 47812 457812 47824
rect 457864 47812 457870 47864
rect 475378 47852 475384 47864
rect 458376 47824 475384 47852
rect 8294 47744 8300 47796
rect 8352 47784 8358 47796
rect 22186 47784 22192 47796
rect 8352 47756 22192 47784
rect 8352 47744 8358 47756
rect 22186 47744 22192 47756
rect 22244 47744 22250 47796
rect 23474 47744 23480 47796
rect 23532 47784 23538 47796
rect 36078 47784 36084 47796
rect 23532 47756 36084 47784
rect 23532 47744 23538 47756
rect 36078 47744 36084 47756
rect 36136 47744 36142 47796
rect 46934 47744 46940 47796
rect 46992 47784 46998 47796
rect 57974 47784 57980 47796
rect 46992 47756 57980 47784
rect 46992 47744 46998 47756
rect 57974 47744 57980 47756
rect 58032 47744 58038 47796
rect 60734 47744 60740 47796
rect 60792 47784 60798 47796
rect 69934 47784 69940 47796
rect 60792 47756 69940 47784
rect 60792 47744 60798 47756
rect 69934 47744 69940 47756
rect 69992 47744 69998 47796
rect 70394 47744 70400 47796
rect 70452 47784 70458 47796
rect 80054 47784 80060 47796
rect 70452 47756 80060 47784
rect 70452 47744 70458 47756
rect 80054 47744 80060 47756
rect 80112 47744 80118 47796
rect 86954 47744 86960 47796
rect 87012 47784 87018 47796
rect 95234 47784 95240 47796
rect 87012 47756 95240 47784
rect 87012 47744 87018 47756
rect 95234 47744 95240 47756
rect 95292 47744 95298 47796
rect 99374 47744 99380 47796
rect 99432 47784 99438 47796
rect 106274 47784 106280 47796
rect 99432 47756 106280 47784
rect 99432 47744 99438 47756
rect 106274 47744 106280 47756
rect 106332 47744 106338 47796
rect 107654 47744 107660 47796
rect 107712 47784 107718 47796
rect 113726 47784 113732 47796
rect 107712 47756 113732 47784
rect 107712 47744 107718 47756
rect 113726 47744 113732 47756
rect 113784 47744 113790 47796
rect 114554 47744 114560 47796
rect 114612 47784 114618 47796
rect 120350 47784 120356 47796
rect 114612 47756 120356 47784
rect 114612 47744 114618 47756
rect 120350 47744 120356 47756
rect 120408 47744 120414 47796
rect 121454 47744 121460 47796
rect 121512 47784 121518 47796
rect 126974 47784 126980 47796
rect 121512 47756 126980 47784
rect 121512 47744 121518 47756
rect 126974 47744 126980 47756
rect 127032 47744 127038 47796
rect 136634 47744 136640 47796
rect 136692 47784 136698 47796
rect 141142 47784 141148 47796
rect 136692 47756 141148 47784
rect 136692 47744 136698 47756
rect 141142 47744 141148 47756
rect 141200 47744 141206 47796
rect 146294 47744 146300 47796
rect 146352 47784 146358 47796
rect 149974 47784 149980 47796
rect 146352 47756 149980 47784
rect 146352 47744 146358 47756
rect 149974 47744 149980 47756
rect 150032 47744 150038 47796
rect 173894 47744 173900 47796
rect 173952 47784 173958 47796
rect 175274 47784 175280 47796
rect 173952 47756 175280 47784
rect 173952 47744 173958 47756
rect 175274 47744 175280 47756
rect 175332 47744 175338 47796
rect 377306 47744 377312 47796
rect 377364 47784 377370 47796
rect 390738 47784 390744 47796
rect 377364 47756 390744 47784
rect 377364 47744 377370 47756
rect 390738 47744 390744 47756
rect 390796 47744 390802 47796
rect 400122 47744 400128 47796
rect 400180 47784 400186 47796
rect 415578 47784 415584 47796
rect 400180 47756 415584 47784
rect 400180 47744 400186 47756
rect 415578 47744 415584 47756
rect 415636 47744 415642 47796
rect 437382 47744 437388 47796
rect 437440 47784 437446 47796
rect 451734 47784 451740 47796
rect 437440 47756 451740 47784
rect 437440 47744 437446 47756
rect 451734 47744 451740 47756
rect 451792 47744 451798 47796
rect 451826 47744 451832 47796
rect 451884 47784 451890 47796
rect 453298 47784 453304 47796
rect 451884 47756 453304 47784
rect 451884 47744 451890 47756
rect 453298 47744 453304 47756
rect 453356 47744 453362 47796
rect 456242 47744 456248 47796
rect 456300 47784 456306 47796
rect 458376 47784 458404 47824
rect 475378 47812 475384 47824
rect 475436 47812 475442 47864
rect 481450 47812 481456 47864
rect 481508 47852 481514 47864
rect 486418 47852 486424 47864
rect 481508 47824 486424 47852
rect 481508 47812 481514 47824
rect 486418 47812 486424 47824
rect 486476 47812 486482 47864
rect 489886 47852 489914 47892
rect 492306 47880 492312 47932
rect 492364 47920 492370 47932
rect 514846 47920 514852 47932
rect 492364 47892 514852 47920
rect 492364 47880 492370 47892
rect 514846 47880 514852 47892
rect 514904 47880 514910 47932
rect 517422 47880 517428 47932
rect 517480 47920 517486 47932
rect 542354 47920 542360 47932
rect 517480 47892 542360 47920
rect 517480 47880 517486 47892
rect 542354 47880 542360 47892
rect 542412 47880 542418 47932
rect 543642 47880 543648 47932
rect 543700 47920 543706 47932
rect 548150 47920 548156 47932
rect 543700 47892 548156 47920
rect 543700 47880 543706 47892
rect 548150 47880 548156 47892
rect 548208 47880 548214 47932
rect 548242 47880 548248 47932
rect 548300 47920 548306 47932
rect 548300 47892 552612 47920
rect 548300 47880 548306 47892
rect 505094 47852 505100 47864
rect 489886 47824 505100 47852
rect 505094 47812 505100 47824
rect 505152 47812 505158 47864
rect 525886 47812 525892 47864
rect 525944 47852 525950 47864
rect 526806 47852 526812 47864
rect 525944 47824 526812 47852
rect 525944 47812 525950 47824
rect 526806 47812 526812 47824
rect 526864 47812 526870 47864
rect 528526 47824 547874 47852
rect 456300 47756 458404 47784
rect 456300 47744 456306 47756
rect 459462 47744 459468 47796
rect 459520 47784 459526 47796
rect 480254 47784 480260 47796
rect 459520 47756 480260 47784
rect 459520 47744 459526 47756
rect 480254 47744 480260 47756
rect 480312 47744 480318 47796
rect 485682 47744 485688 47796
rect 485740 47784 485746 47796
rect 507854 47784 507860 47796
rect 485740 47756 507860 47784
rect 485740 47744 485746 47756
rect 507854 47744 507860 47756
rect 507912 47744 507918 47796
rect 525242 47744 525248 47796
rect 525300 47784 525306 47796
rect 528526 47784 528554 47824
rect 525300 47756 528554 47784
rect 547846 47784 547874 47824
rect 549162 47812 549168 47864
rect 549220 47852 549226 47864
rect 551278 47852 551284 47864
rect 549220 47824 551284 47852
rect 549220 47812 549226 47824
rect 551278 47812 551284 47824
rect 551336 47812 551342 47864
rect 550634 47784 550640 47796
rect 547846 47756 550640 47784
rect 525300 47744 525306 47756
rect 550634 47744 550640 47756
rect 550692 47744 550698 47796
rect 552584 47784 552612 47892
rect 552658 47812 552664 47864
rect 552716 47852 552722 47864
rect 560938 47852 560944 47864
rect 552716 47824 560944 47852
rect 552716 47812 552722 47824
rect 560938 47812 560944 47824
rect 560996 47812 561002 47864
rect 566458 47784 566464 47796
rect 552584 47756 566464 47784
rect 566458 47744 566464 47756
rect 566516 47744 566522 47796
rect 6914 47676 6920 47728
rect 6972 47716 6978 47728
rect 20714 47716 20720 47728
rect 6972 47688 20720 47716
rect 6972 47676 6978 47688
rect 20714 47676 20720 47688
rect 20772 47676 20778 47728
rect 27614 47676 27620 47728
rect 27672 47716 27678 47728
rect 40310 47716 40316 47728
rect 27672 47688 40316 47716
rect 27672 47676 27678 47688
rect 40310 47676 40316 47688
rect 40368 47676 40374 47728
rect 48406 47676 48412 47728
rect 48464 47716 48470 47728
rect 59446 47716 59452 47728
rect 48464 47688 59452 47716
rect 48464 47676 48470 47688
rect 59446 47676 59452 47688
rect 59504 47676 59510 47728
rect 62114 47676 62120 47728
rect 62172 47716 62178 47728
rect 72142 47716 72148 47728
rect 62172 47688 72148 47716
rect 62172 47676 62178 47688
rect 72142 47676 72148 47688
rect 72200 47676 72206 47728
rect 75914 47676 75920 47728
rect 75972 47716 75978 47728
rect 84286 47716 84292 47728
rect 75972 47688 84292 47716
rect 75972 47676 75978 47688
rect 84286 47676 84292 47688
rect 84344 47676 84350 47728
rect 88334 47676 88340 47728
rect 88392 47716 88398 47728
rect 96706 47716 96712 47728
rect 88392 47688 96712 47716
rect 88392 47676 88398 47688
rect 96706 47676 96712 47688
rect 96764 47676 96770 47728
rect 102318 47676 102324 47728
rect 102376 47716 102382 47728
rect 109310 47716 109316 47728
rect 102376 47688 109316 47716
rect 102376 47676 102382 47688
rect 109310 47676 109316 47688
rect 109368 47676 109374 47728
rect 110598 47676 110604 47728
rect 110656 47716 110662 47728
rect 115934 47716 115940 47728
rect 110656 47688 115940 47716
rect 110656 47676 110662 47688
rect 115934 47676 115940 47688
rect 115992 47676 115998 47728
rect 124306 47676 124312 47728
rect 124364 47716 124370 47728
rect 129182 47716 129188 47728
rect 124364 47688 129188 47716
rect 124364 47676 124370 47688
rect 129182 47676 129188 47688
rect 129240 47676 129246 47728
rect 132586 47676 132592 47728
rect 132644 47716 132650 47728
rect 136726 47716 136732 47728
rect 132644 47688 136732 47716
rect 132644 47676 132650 47688
rect 136726 47676 136732 47688
rect 136784 47676 136790 47728
rect 151906 47676 151912 47728
rect 151964 47716 151970 47728
rect 154574 47716 154580 47728
rect 151964 47688 154580 47716
rect 151964 47676 151970 47688
rect 154574 47676 154580 47688
rect 154632 47676 154638 47728
rect 362862 47676 362868 47728
rect 362920 47716 362926 47728
rect 375374 47716 375380 47728
rect 362920 47688 375380 47716
rect 362920 47676 362926 47688
rect 375374 47676 375380 47688
rect 375432 47676 375438 47728
rect 380618 47676 380624 47728
rect 380676 47716 380682 47728
rect 394694 47716 394700 47728
rect 380676 47688 394700 47716
rect 380676 47676 380682 47688
rect 394694 47676 394700 47688
rect 394752 47676 394758 47728
rect 396994 47676 397000 47728
rect 397052 47716 397058 47728
rect 412634 47716 412640 47728
rect 397052 47688 412640 47716
rect 397052 47676 397058 47688
rect 412634 47676 412640 47688
rect 412692 47676 412698 47728
rect 426342 47676 426348 47728
rect 426400 47716 426406 47728
rect 444374 47716 444380 47728
rect 426400 47688 444380 47716
rect 426400 47676 426406 47688
rect 444374 47676 444380 47688
rect 444432 47676 444438 47728
rect 449618 47676 449624 47728
rect 449676 47716 449682 47728
rect 469214 47716 469220 47728
rect 449676 47688 469220 47716
rect 449676 47676 449682 47688
rect 469214 47676 469220 47688
rect 469272 47676 469278 47728
rect 472618 47676 472624 47728
rect 472676 47716 472682 47728
rect 494054 47716 494060 47728
rect 472676 47688 494060 47716
rect 472676 47676 472682 47688
rect 494054 47676 494060 47688
rect 494112 47676 494118 47728
rect 495250 47676 495256 47728
rect 495308 47716 495314 47728
rect 518894 47716 518900 47728
rect 495308 47688 518900 47716
rect 495308 47676 495314 47688
rect 518894 47676 518900 47688
rect 518952 47676 518958 47728
rect 536098 47676 536104 47728
rect 536156 47716 536162 47728
rect 563054 47716 563060 47728
rect 536156 47688 563060 47716
rect 536156 47676 536162 47688
rect 563054 47676 563060 47688
rect 563112 47676 563118 47728
rect 5534 47608 5540 47660
rect 5592 47648 5598 47660
rect 19518 47648 19524 47660
rect 5592 47620 19524 47648
rect 5592 47608 5598 47620
rect 19518 47608 19524 47620
rect 19576 47608 19582 47660
rect 28994 47608 29000 47660
rect 29052 47648 29058 47660
rect 41414 47648 41420 47660
rect 29052 47620 41420 47648
rect 29052 47608 29058 47620
rect 41414 47608 41420 47620
rect 41472 47608 41478 47660
rect 42794 47608 42800 47660
rect 42852 47648 42858 47660
rect 53926 47648 53932 47660
rect 42852 47620 53932 47648
rect 42852 47608 42858 47620
rect 53926 47608 53932 47620
rect 53984 47608 53990 47660
rect 57974 47608 57980 47660
rect 58032 47648 58038 47660
rect 67726 47648 67732 47660
rect 58032 47620 67732 47648
rect 58032 47608 58038 47620
rect 67726 47608 67732 47620
rect 67784 47608 67790 47660
rect 69014 47608 69020 47660
rect 69072 47648 69078 47660
rect 78858 47648 78864 47660
rect 69072 47620 78864 47648
rect 69072 47608 69078 47620
rect 78858 47608 78864 47620
rect 78916 47608 78922 47660
rect 81434 47608 81440 47660
rect 81492 47648 81498 47660
rect 89714 47648 89720 47660
rect 81492 47620 89720 47648
rect 81492 47608 81498 47620
rect 89714 47608 89720 47620
rect 89772 47608 89778 47660
rect 95234 47608 95240 47660
rect 95292 47648 95298 47660
rect 102870 47648 102876 47660
rect 95292 47620 102876 47648
rect 95292 47608 95298 47620
rect 102870 47608 102876 47620
rect 102928 47608 102934 47660
rect 106274 47608 106280 47660
rect 106332 47648 106338 47660
rect 112622 47648 112628 47660
rect 106332 47620 112628 47648
rect 106332 47608 106338 47620
rect 112622 47608 112628 47620
rect 112680 47608 112686 47660
rect 131206 47608 131212 47660
rect 131264 47648 131270 47660
rect 135622 47648 135628 47660
rect 131264 47620 135628 47648
rect 131264 47608 131270 47620
rect 135622 47608 135628 47620
rect 135680 47608 135686 47660
rect 137278 47608 137284 47660
rect 137336 47648 137342 47660
rect 140038 47648 140044 47660
rect 137336 47620 140044 47648
rect 137336 47608 137342 47620
rect 140038 47608 140044 47620
rect 140096 47608 140102 47660
rect 147766 47608 147772 47660
rect 147824 47648 147830 47660
rect 151078 47648 151084 47660
rect 147824 47620 151084 47648
rect 147824 47608 147830 47620
rect 151078 47608 151084 47620
rect 151136 47608 151142 47660
rect 158806 47608 158812 47660
rect 158864 47648 158870 47660
rect 160830 47648 160836 47660
rect 158864 47620 160836 47648
rect 158864 47608 158870 47620
rect 160830 47608 160836 47620
rect 160888 47608 160894 47660
rect 162946 47608 162952 47660
rect 163004 47648 163010 47660
rect 165614 47648 165620 47660
rect 163004 47620 165620 47648
rect 163004 47608 163010 47620
rect 165614 47608 165620 47620
rect 165672 47608 165678 47660
rect 168374 47608 168380 47660
rect 168432 47648 168438 47660
rect 169754 47648 169760 47660
rect 168432 47620 169760 47648
rect 168432 47608 168438 47620
rect 169754 47608 169760 47620
rect 169812 47608 169818 47660
rect 234614 47608 234620 47660
rect 234672 47648 234678 47660
rect 237374 47648 237380 47660
rect 234672 47620 237380 47648
rect 234672 47608 234678 47620
rect 237374 47608 237380 47620
rect 237432 47608 237438 47660
rect 239950 47608 239956 47660
rect 240008 47648 240014 47660
rect 240778 47648 240784 47660
rect 240008 47620 240784 47648
rect 240008 47608 240014 47620
rect 240778 47608 240784 47620
rect 240836 47608 240842 47660
rect 243722 47608 243728 47660
rect 243780 47648 243786 47660
rect 246298 47648 246304 47660
rect 243780 47620 246304 47648
rect 243780 47608 243786 47620
rect 246298 47608 246304 47620
rect 246356 47608 246362 47660
rect 350626 47608 350632 47660
rect 350684 47648 350690 47660
rect 362218 47648 362224 47660
rect 350684 47620 362224 47648
rect 350684 47608 350690 47620
rect 362218 47608 362224 47620
rect 362276 47608 362282 47660
rect 367094 47608 367100 47660
rect 367152 47648 367158 47660
rect 380894 47648 380900 47660
rect 367152 47620 380900 47648
rect 367152 47608 367158 47620
rect 380894 47608 380900 47620
rect 380952 47608 380958 47660
rect 383470 47608 383476 47660
rect 383528 47648 383534 47660
rect 399018 47648 399024 47660
rect 383528 47620 399024 47648
rect 383528 47608 383534 47620
rect 399018 47608 399024 47620
rect 399076 47608 399082 47660
rect 403618 47608 403624 47660
rect 403676 47648 403682 47660
rect 419534 47648 419540 47660
rect 403676 47620 419540 47648
rect 403676 47608 403682 47620
rect 419534 47608 419540 47620
rect 419592 47608 419598 47660
rect 420730 47608 420736 47660
rect 420788 47648 420794 47660
rect 438118 47648 438124 47660
rect 420788 47620 438124 47648
rect 420788 47608 420794 47620
rect 438118 47608 438124 47620
rect 438176 47608 438182 47660
rect 442902 47608 442908 47660
rect 442960 47648 442966 47660
rect 462314 47648 462320 47660
rect 442960 47620 462320 47648
rect 442960 47608 442966 47620
rect 462314 47608 462320 47620
rect 462372 47608 462378 47660
rect 468202 47608 468208 47660
rect 468260 47648 468266 47660
rect 490006 47648 490012 47660
rect 468260 47620 490012 47648
rect 468260 47608 468266 47620
rect 490006 47608 490012 47620
rect 490064 47608 490070 47660
rect 498930 47608 498936 47660
rect 498988 47648 498994 47660
rect 523218 47648 523224 47660
rect 498988 47620 523224 47648
rect 498988 47608 498994 47620
rect 523218 47608 523224 47620
rect 523276 47608 523282 47660
rect 528278 47608 528284 47660
rect 528336 47648 528342 47660
rect 554774 47648 554780 47660
rect 528336 47620 554780 47648
rect 528336 47608 528342 47620
rect 554774 47608 554780 47620
rect 554832 47608 554838 47660
rect 4154 47540 4160 47592
rect 4212 47580 4218 47592
rect 18414 47580 18420 47592
rect 4212 47552 18420 47580
rect 4212 47540 4218 47552
rect 18414 47540 18420 47552
rect 18472 47540 18478 47592
rect 20714 47540 20720 47592
rect 20772 47580 20778 47592
rect 33870 47580 33876 47592
rect 20772 47552 33876 47580
rect 20772 47540 20778 47552
rect 33870 47540 33876 47552
rect 33928 47540 33934 47592
rect 35894 47540 35900 47592
rect 35952 47580 35958 47592
rect 48314 47580 48320 47592
rect 35952 47552 48320 47580
rect 35952 47540 35958 47552
rect 48314 47540 48320 47552
rect 48372 47540 48378 47592
rect 52454 47540 52460 47592
rect 52512 47580 52518 47592
rect 63494 47580 63500 47592
rect 52512 47552 63500 47580
rect 52512 47540 52518 47552
rect 63494 47540 63500 47552
rect 63552 47540 63558 47592
rect 64874 47540 64880 47592
rect 64932 47580 64938 47592
rect 74534 47580 74540 47592
rect 64932 47552 74540 47580
rect 64932 47540 64938 47552
rect 74534 47540 74540 47552
rect 74592 47540 74598 47592
rect 75178 47540 75184 47592
rect 75236 47580 75242 47592
rect 82078 47580 82084 47592
rect 75236 47552 82084 47580
rect 75236 47540 75242 47552
rect 82078 47540 82084 47552
rect 82136 47540 82142 47592
rect 82814 47540 82820 47592
rect 82872 47580 82878 47592
rect 91186 47580 91192 47592
rect 82872 47552 91192 47580
rect 82872 47540 82878 47552
rect 91186 47540 91192 47552
rect 91244 47540 91250 47592
rect 93946 47540 93952 47592
rect 94004 47580 94010 47592
rect 101766 47580 101772 47592
rect 94004 47552 101772 47580
rect 94004 47540 94010 47552
rect 101766 47540 101772 47552
rect 101824 47540 101830 47592
rect 110506 47540 110512 47592
rect 110564 47580 110570 47592
rect 117314 47580 117320 47592
rect 110564 47552 117320 47580
rect 110564 47540 110570 47552
rect 117314 47540 117320 47552
rect 117372 47540 117378 47592
rect 122834 47540 122840 47592
rect 122892 47580 122898 47592
rect 128446 47580 128452 47592
rect 122892 47552 128452 47580
rect 122892 47540 122898 47552
rect 128446 47540 128452 47552
rect 128504 47540 128510 47592
rect 143626 47540 143632 47592
rect 143684 47580 143690 47592
rect 147858 47580 147864 47592
rect 143684 47552 147864 47580
rect 143684 47540 143690 47552
rect 147858 47540 147864 47552
rect 147916 47540 147922 47592
rect 154574 47540 154580 47592
rect 154632 47580 154638 47592
rect 157518 47580 157524 47592
rect 154632 47552 157524 47580
rect 154632 47540 154638 47552
rect 157518 47540 157524 47552
rect 157576 47540 157582 47592
rect 265618 47540 265624 47592
rect 265676 47580 265682 47592
rect 270494 47580 270500 47592
rect 265676 47552 270500 47580
rect 265676 47540 265682 47552
rect 270494 47540 270500 47552
rect 270552 47540 270558 47592
rect 293862 47540 293868 47592
rect 293920 47580 293926 47592
rect 300118 47580 300124 47592
rect 293920 47552 300124 47580
rect 293920 47540 293926 47552
rect 300118 47540 300124 47552
rect 300176 47540 300182 47592
rect 347682 47540 347688 47592
rect 347740 47580 347746 47592
rect 358078 47580 358084 47592
rect 347740 47552 358084 47580
rect 347740 47540 347746 47552
rect 358078 47540 358084 47552
rect 358136 47540 358142 47592
rect 373810 47540 373816 47592
rect 373868 47580 373874 47592
rect 387794 47580 387800 47592
rect 373868 47552 387800 47580
rect 373868 47540 373874 47552
rect 387794 47540 387800 47552
rect 387852 47540 387858 47592
rect 390370 47540 390376 47592
rect 390428 47580 390434 47592
rect 405734 47580 405740 47592
rect 390428 47552 405740 47580
rect 390428 47540 390434 47552
rect 405734 47540 405740 47552
rect 405792 47540 405798 47592
rect 406930 47540 406936 47592
rect 406988 47580 406994 47592
rect 423858 47580 423864 47592
rect 406988 47552 423864 47580
rect 406988 47540 406994 47552
rect 423858 47540 423864 47552
rect 423916 47540 423922 47592
rect 429930 47540 429936 47592
rect 429988 47580 429994 47592
rect 448606 47580 448612 47592
rect 429988 47552 448612 47580
rect 429988 47540 429994 47552
rect 448606 47540 448612 47552
rect 448664 47540 448670 47592
rect 451734 47540 451740 47592
rect 451792 47580 451798 47592
rect 457070 47580 457076 47592
rect 451792 47552 457076 47580
rect 451792 47540 451798 47552
rect 457070 47540 457076 47552
rect 457128 47540 457134 47592
rect 473538 47580 473544 47592
rect 460906 47552 473544 47580
rect 9674 47472 9680 47524
rect 9732 47512 9738 47524
rect 22830 47512 22836 47524
rect 9732 47484 22836 47512
rect 9732 47472 9738 47484
rect 22830 47472 22836 47484
rect 22888 47472 22894 47524
rect 26234 47472 26240 47524
rect 26292 47512 26298 47524
rect 38102 47512 38108 47524
rect 26292 47484 38108 47512
rect 26292 47472 26298 47484
rect 38102 47472 38108 47484
rect 38160 47472 38166 47524
rect 49694 47472 49700 47524
rect 49752 47512 49758 47524
rect 60182 47512 60188 47524
rect 49752 47484 60188 47512
rect 49752 47472 49758 47484
rect 60182 47472 60188 47484
rect 60240 47472 60246 47524
rect 84286 47472 84292 47524
rect 84344 47512 84350 47524
rect 91830 47512 91836 47524
rect 84344 47484 91836 47512
rect 84344 47472 84350 47484
rect 91830 47472 91836 47484
rect 91888 47472 91894 47524
rect 142154 47472 142160 47524
rect 142212 47512 142218 47524
rect 145558 47512 145564 47524
rect 142212 47484 145564 47512
rect 142212 47472 142218 47484
rect 145558 47472 145564 47484
rect 145616 47472 145622 47524
rect 156046 47472 156052 47524
rect 156104 47512 156110 47524
rect 158714 47512 158720 47524
rect 156104 47484 158720 47512
rect 156104 47472 156110 47484
rect 158714 47472 158720 47484
rect 158772 47472 158778 47524
rect 427722 47472 427728 47524
rect 427780 47512 427786 47524
rect 439498 47512 439504 47524
rect 427780 47484 439504 47512
rect 427780 47472 427786 47484
rect 439498 47472 439504 47484
rect 439556 47472 439562 47524
rect 452470 47472 452476 47524
rect 452528 47512 452534 47524
rect 460906 47512 460934 47552
rect 473538 47540 473544 47552
rect 473596 47540 473602 47592
rect 475930 47540 475936 47592
rect 475988 47580 475994 47592
rect 498194 47580 498200 47592
rect 475988 47552 498200 47580
rect 475988 47540 475994 47552
rect 498194 47540 498200 47552
rect 498252 47540 498258 47592
rect 502242 47540 502248 47592
rect 502300 47580 502306 47592
rect 525794 47580 525800 47592
rect 502300 47552 525800 47580
rect 502300 47540 502306 47552
rect 525794 47540 525800 47552
rect 525852 47540 525858 47592
rect 534994 47540 535000 47592
rect 535052 47580 535058 47592
rect 561674 47580 561680 47592
rect 535052 47552 561680 47580
rect 535052 47540 535058 47552
rect 561674 47540 561680 47552
rect 561732 47540 561738 47592
rect 452528 47484 460934 47512
rect 452528 47472 452534 47484
rect 481266 47472 481272 47524
rect 481324 47512 481330 47524
rect 487154 47512 487160 47524
rect 481324 47484 487160 47512
rect 481324 47472 481330 47484
rect 487154 47472 487160 47484
rect 487212 47472 487218 47524
rect 521470 47472 521476 47524
rect 521528 47512 521534 47524
rect 548058 47512 548064 47524
rect 521528 47484 548064 47512
rect 521528 47472 521534 47484
rect 548058 47472 548064 47484
rect 548116 47472 548122 47524
rect 548150 47472 548156 47524
rect 548208 47512 548214 47524
rect 556798 47512 556804 47524
rect 548208 47484 556804 47512
rect 548208 47472 548214 47484
rect 556798 47472 556804 47484
rect 556856 47472 556862 47524
rect 17954 47404 17960 47456
rect 18012 47444 18018 47456
rect 30558 47444 30564 47456
rect 18012 47416 30564 47444
rect 18012 47404 18018 47416
rect 30558 47404 30564 47416
rect 30616 47404 30622 47456
rect 34514 47404 34520 47456
rect 34572 47444 34578 47456
rect 45830 47444 45836 47456
rect 34572 47416 45836 47444
rect 34572 47404 34578 47416
rect 45830 47404 45836 47416
rect 45888 47404 45894 47456
rect 74534 47404 74540 47456
rect 74592 47444 74598 47456
rect 83182 47444 83188 47456
rect 74592 47416 83188 47444
rect 74592 47404 74598 47416
rect 83182 47404 83188 47416
rect 83240 47404 83246 47456
rect 207474 47404 207480 47456
rect 207532 47444 207538 47456
rect 208394 47444 208400 47456
rect 207532 47416 208400 47444
rect 207532 47404 207538 47416
rect 208394 47404 208400 47416
rect 208452 47404 208458 47456
rect 13906 47336 13912 47388
rect 13964 47376 13970 47388
rect 27246 47376 27252 47388
rect 13964 47348 27252 47376
rect 13964 47336 13970 47348
rect 27246 47336 27252 47348
rect 27304 47336 27310 47388
rect 37274 47336 37280 47388
rect 37332 47376 37338 47388
rect 49142 47376 49148 47388
rect 37332 47348 49148 47376
rect 37332 47336 37338 47348
rect 49142 47336 49148 47348
rect 49200 47336 49206 47388
rect 135438 47336 135444 47388
rect 135496 47376 135502 47388
rect 138934 47376 138940 47388
rect 135496 47348 138940 47376
rect 135496 47336 135502 47348
rect 138934 47336 138940 47348
rect 138992 47336 138998 47388
rect 165614 47336 165620 47388
rect 165672 47376 165678 47388
rect 167454 47376 167460 47388
rect 165672 47348 167460 47376
rect 165672 47336 165678 47348
rect 167454 47336 167460 47348
rect 167512 47336 167518 47388
rect 519722 47336 519728 47388
rect 519780 47376 519786 47388
rect 522298 47376 522304 47388
rect 519780 47348 522304 47376
rect 519780 47336 519786 47348
rect 522298 47336 522304 47348
rect 522356 47336 522362 47388
rect 551554 47336 551560 47388
rect 551612 47376 551618 47388
rect 558178 47376 558184 47388
rect 551612 47348 558184 47376
rect 551612 47336 551618 47348
rect 558178 47336 558184 47348
rect 558236 47336 558242 47388
rect 27706 47268 27712 47320
rect 27764 47308 27770 47320
rect 39206 47308 39212 47320
rect 27764 47280 39212 47308
rect 27764 47268 27770 47280
rect 39206 47268 39212 47280
rect 39264 47268 39270 47320
rect 44266 47268 44272 47320
rect 44324 47308 44330 47320
rect 54662 47308 54668 47320
rect 44324 47280 54668 47308
rect 44324 47268 44330 47280
rect 54662 47268 54668 47280
rect 54720 47268 54726 47320
rect 85574 47268 85580 47320
rect 85632 47308 85638 47320
rect 92934 47308 92940 47320
rect 85632 47280 92940 47308
rect 85632 47268 85638 47280
rect 92934 47268 92940 47280
rect 92992 47268 92998 47320
rect 93854 47268 93860 47320
rect 93912 47308 93918 47320
rect 100754 47308 100760 47320
rect 93912 47280 100760 47308
rect 93912 47268 93918 47280
rect 100754 47268 100760 47280
rect 100812 47268 100818 47320
rect 237098 47268 237104 47320
rect 237156 47308 237162 47320
rect 240134 47308 240140 47320
rect 237156 47280 240140 47308
rect 237156 47268 237162 47280
rect 240134 47268 240140 47280
rect 240192 47268 240198 47320
rect 522942 47268 522948 47320
rect 523000 47308 523006 47320
rect 529198 47308 529204 47320
rect 523000 47280 529204 47308
rect 523000 47268 523006 47280
rect 529198 47268 529204 47280
rect 529256 47268 529262 47320
rect 25498 47200 25504 47252
rect 25556 47240 25562 47252
rect 32766 47240 32772 47252
rect 25556 47212 32772 47240
rect 25556 47200 25562 47212
rect 32766 47200 32772 47212
rect 32824 47200 32830 47252
rect 124858 47200 124864 47252
rect 124916 47240 124922 47252
rect 125870 47240 125876 47252
rect 124916 47212 125876 47240
rect 124916 47200 124922 47212
rect 125870 47200 125876 47212
rect 125928 47200 125934 47252
rect 172514 47200 172520 47252
rect 172572 47240 172578 47252
rect 174078 47240 174084 47252
rect 172572 47212 174084 47240
rect 172572 47200 172578 47212
rect 174078 47200 174084 47212
rect 174136 47200 174142 47252
rect 117314 47064 117320 47116
rect 117372 47104 117378 47116
rect 122926 47104 122932 47116
rect 117372 47076 122932 47104
rect 117372 47064 117378 47076
rect 122926 47064 122932 47076
rect 122984 47064 122990 47116
rect 118786 46996 118792 47048
rect 118844 47036 118850 47048
rect 124766 47036 124772 47048
rect 118844 47008 124772 47036
rect 118844 46996 118850 47008
rect 124766 46996 124772 47008
rect 124824 46996 124830 47048
rect 130378 46996 130384 47048
rect 130436 47036 130442 47048
rect 133414 47036 133420 47048
rect 130436 47008 133420 47036
rect 130436 46996 130442 47008
rect 133414 46996 133420 47008
rect 133472 46996 133478 47048
rect 139486 46996 139492 47048
rect 139544 47036 139550 47048
rect 143534 47036 143540 47048
rect 139544 47008 143540 47036
rect 139544 46996 139550 47008
rect 143534 46996 143540 47008
rect 143592 46996 143598 47048
rect 150526 46996 150532 47048
rect 150584 47036 150590 47048
rect 153286 47036 153292 47048
rect 150584 47008 153292 47036
rect 150584 46996 150590 47008
rect 153286 46996 153292 47008
rect 153344 46996 153350 47048
rect 160094 46996 160100 47048
rect 160152 47036 160158 47048
rect 163038 47036 163044 47048
rect 160152 47008 163044 47036
rect 160152 46996 160158 47008
rect 163038 46996 163044 47008
rect 163096 46996 163102 47048
rect 77294 46928 77300 46980
rect 77352 46968 77358 46980
rect 86310 46968 86316 46980
rect 77352 46940 86316 46968
rect 77352 46928 77358 46940
rect 86310 46928 86316 46940
rect 86368 46928 86374 46980
rect 118878 46928 118884 46980
rect 118936 46968 118942 46980
rect 123662 46968 123668 46980
rect 118936 46940 123668 46968
rect 118936 46928 118942 46940
rect 123662 46928 123668 46940
rect 123720 46928 123726 46980
rect 140866 46928 140872 46980
rect 140924 46968 140930 46980
rect 144454 46968 144460 46980
rect 140924 46940 144460 46968
rect 140924 46928 140930 46940
rect 144454 46928 144460 46940
rect 144512 46928 144518 46980
rect 149238 46928 149244 46980
rect 149296 46968 149302 46980
rect 152182 46968 152188 46980
rect 149296 46940 152188 46968
rect 149296 46928 149302 46940
rect 152182 46928 152188 46940
rect 152240 46928 152246 46980
rect 160278 46928 160284 46980
rect 160336 46968 160342 46980
rect 161934 46968 161940 46980
rect 160336 46940 161940 46968
rect 160336 46928 160342 46940
rect 161934 46928 161940 46940
rect 161992 46928 161998 46980
rect 169754 46928 169760 46980
rect 169812 46968 169818 46980
rect 171870 46968 171876 46980
rect 169812 46940 171876 46968
rect 169812 46928 169818 46940
rect 171870 46928 171876 46940
rect 171928 46928 171934 46980
rect 179414 46928 179420 46980
rect 179472 46968 179478 46980
rect 180794 46968 180800 46980
rect 179472 46940 180800 46968
rect 179472 46928 179478 46940
rect 180794 46928 180800 46940
rect 180852 46928 180858 46980
rect 219342 46928 219348 46980
rect 219400 46968 219406 46980
rect 220078 46968 220084 46980
rect 219400 46940 220084 46968
rect 219400 46928 219406 46940
rect 220078 46928 220084 46940
rect 220136 46928 220142 46980
rect 362034 46928 362040 46980
rect 362092 46968 362098 46980
rect 366358 46968 366364 46980
rect 362092 46940 366364 46968
rect 362092 46928 362098 46940
rect 366358 46928 366364 46940
rect 366416 46928 366422 46980
rect 487890 46928 487896 46980
rect 487948 46968 487954 46980
rect 490558 46968 490564 46980
rect 487948 46940 490564 46968
rect 487948 46928 487954 46940
rect 490558 46928 490564 46940
rect 490616 46928 490622 46980
rect 223574 46452 223580 46504
rect 223632 46492 223638 46504
rect 224494 46492 224500 46504
rect 223632 46464 224500 46492
rect 223632 46452 223638 46464
rect 224494 46452 224500 46464
rect 224552 46452 224558 46504
rect 160094 11704 160100 11756
rect 160152 11744 160158 11756
rect 161290 11744 161296 11756
rect 160152 11716 161296 11744
rect 160152 11704 160158 11716
rect 161290 11704 161296 11716
rect 161348 11704 161354 11756
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 516134 5448 516140 5500
rect 516192 5488 516198 5500
rect 541986 5488 541992 5500
rect 516192 5460 541992 5488
rect 516192 5448 516198 5460
rect 541986 5448 541992 5460
rect 542044 5448 542050 5500
rect 525978 5380 525984 5432
rect 526036 5420 526042 5432
rect 552658 5420 552664 5432
rect 526036 5392 552664 5420
rect 526036 5380 526042 5392
rect 552658 5380 552664 5392
rect 552716 5380 552722 5432
rect 517514 5312 517520 5364
rect 517572 5352 517578 5364
rect 544378 5352 544384 5364
rect 517572 5324 544384 5352
rect 517572 5312 517578 5324
rect 544378 5312 544384 5324
rect 544436 5312 544442 5364
rect 531314 5244 531320 5296
rect 531372 5284 531378 5296
rect 558546 5284 558552 5296
rect 531372 5256 558552 5284
rect 531372 5244 531378 5256
rect 558546 5244 558552 5256
rect 558604 5244 558610 5296
rect 473354 5176 473360 5228
rect 473412 5216 473418 5228
rect 495894 5216 495900 5228
rect 473412 5188 495900 5216
rect 473412 5176 473418 5188
rect 495894 5176 495900 5188
rect 495952 5176 495958 5228
rect 505186 5176 505192 5228
rect 505244 5216 505250 5228
rect 530118 5216 530124 5228
rect 505244 5188 530124 5216
rect 505244 5176 505250 5188
rect 530118 5176 530124 5188
rect 530176 5176 530182 5228
rect 531498 5176 531504 5228
rect 531556 5216 531562 5228
rect 559742 5216 559748 5228
rect 531556 5188 559748 5216
rect 531556 5176 531562 5188
rect 559742 5176 559748 5188
rect 559800 5176 559806 5228
rect 469306 5108 469312 5160
rect 469364 5148 469370 5160
rect 492306 5148 492312 5160
rect 469364 5120 492312 5148
rect 469364 5108 469370 5120
rect 492306 5108 492312 5120
rect 492364 5108 492370 5160
rect 509234 5108 509240 5160
rect 509292 5148 509298 5160
rect 534902 5148 534908 5160
rect 509292 5120 534908 5148
rect 509292 5108 509298 5120
rect 534902 5108 534908 5120
rect 534960 5108 534966 5160
rect 542446 5108 542452 5160
rect 542504 5148 542510 5160
rect 570322 5148 570328 5160
rect 542504 5120 570328 5148
rect 542504 5108 542510 5120
rect 570322 5108 570328 5120
rect 570380 5108 570386 5160
rect 488534 5040 488540 5092
rect 488592 5080 488598 5092
rect 513558 5080 513564 5092
rect 488592 5052 513564 5080
rect 488592 5040 488598 5052
rect 513558 5040 513564 5052
rect 513616 5040 513622 5092
rect 528554 5040 528560 5092
rect 528612 5080 528618 5092
rect 556154 5080 556160 5092
rect 528612 5052 556160 5080
rect 528612 5040 528618 5052
rect 556154 5040 556160 5052
rect 556212 5040 556218 5092
rect 478874 4972 478880 5024
rect 478932 5012 478938 5024
rect 501782 5012 501788 5024
rect 478932 4984 501788 5012
rect 478932 4972 478938 4984
rect 501782 4972 501788 4984
rect 501840 4972 501846 5024
rect 502334 4972 502340 5024
rect 502392 5012 502398 5024
rect 527818 5012 527824 5024
rect 502392 4984 527824 5012
rect 502392 4972 502398 4984
rect 527818 4972 527824 4984
rect 527876 4972 527882 5024
rect 538214 4972 538220 5024
rect 538272 5012 538278 5024
rect 566826 5012 566832 5024
rect 538272 4984 566832 5012
rect 538272 4972 538278 4984
rect 566826 4972 566832 4984
rect 566884 4972 566890 5024
rect 466454 4904 466460 4956
rect 466512 4944 466518 4956
rect 488810 4944 488816 4956
rect 466512 4916 488816 4944
rect 466512 4904 466518 4916
rect 488810 4904 488816 4916
rect 488868 4904 488874 4956
rect 495434 4904 495440 4956
rect 495492 4944 495498 4956
rect 520734 4944 520740 4956
rect 495492 4916 520740 4944
rect 495492 4904 495498 4916
rect 520734 4904 520740 4916
rect 520792 4904 520798 4956
rect 536834 4904 536840 4956
rect 536892 4944 536898 4956
rect 565630 4944 565636 4956
rect 536892 4916 565636 4944
rect 536892 4904 536898 4916
rect 565630 4904 565636 4916
rect 565688 4904 565694 4956
rect 476114 4836 476120 4888
rect 476172 4876 476178 4888
rect 499390 4876 499396 4888
rect 476172 4848 499396 4876
rect 476172 4836 476178 4848
rect 499390 4836 499396 4848
rect 499448 4836 499454 4888
rect 505278 4836 505284 4888
rect 505336 4876 505342 4888
rect 531314 4876 531320 4888
rect 505336 4848 531320 4876
rect 505336 4836 505342 4848
rect 531314 4836 531320 4848
rect 531372 4836 531378 4888
rect 540974 4836 540980 4888
rect 541032 4876 541038 4888
rect 569126 4876 569132 4888
rect 541032 4848 569132 4876
rect 541032 4836 541038 4848
rect 569126 4836 569132 4848
rect 569184 4836 569190 4888
rect 440326 4768 440332 4820
rect 440384 4808 440390 4820
rect 460382 4808 460388 4820
rect 440384 4780 460388 4808
rect 440384 4768 440390 4780
rect 460382 4768 460388 4780
rect 460440 4768 460446 4820
rect 478966 4768 478972 4820
rect 479024 4808 479030 4820
rect 502978 4808 502984 4820
rect 479024 4780 502984 4808
rect 479024 4768 479030 4780
rect 502978 4768 502984 4780
rect 503036 4768 503042 4820
rect 510706 4768 510712 4820
rect 510764 4808 510770 4820
rect 537202 4808 537208 4820
rect 510764 4780 537208 4808
rect 510764 4768 510770 4780
rect 537202 4768 537208 4780
rect 537260 4768 537266 4820
rect 543734 4768 543740 4820
rect 543792 4808 543798 4820
rect 572714 4808 572720 4820
rect 543792 4780 572720 4808
rect 543792 4768 543798 4780
rect 572714 4768 572720 4780
rect 572772 4768 572778 4820
rect 77386 4088 77392 4140
rect 77444 4128 77450 4140
rect 85758 4128 85764 4140
rect 77444 4100 85764 4128
rect 77444 4088 77450 4100
rect 85758 4088 85764 4100
rect 85816 4088 85822 4140
rect 252554 4088 252560 4140
rect 252612 4128 252618 4140
rect 258258 4128 258264 4140
rect 252612 4100 258264 4128
rect 252612 4088 252618 4100
rect 258258 4088 258264 4100
rect 258316 4088 258322 4140
rect 292574 4088 292580 4140
rect 292632 4128 292638 4140
rect 300762 4128 300768 4140
rect 292632 4100 300768 4128
rect 292632 4088 292638 4100
rect 300762 4088 300768 4100
rect 300820 4088 300826 4140
rect 302234 4088 302240 4140
rect 302292 4128 302298 4140
rect 311434 4128 311440 4140
rect 302292 4100 311440 4128
rect 302292 4088 302298 4100
rect 311434 4088 311440 4100
rect 311492 4088 311498 4140
rect 313274 4088 313280 4140
rect 313332 4128 313338 4140
rect 324406 4128 324412 4140
rect 313332 4100 324412 4128
rect 313332 4088 313338 4100
rect 324406 4088 324412 4100
rect 324464 4088 324470 4140
rect 339494 4088 339500 4140
rect 339552 4128 339558 4140
rect 351638 4128 351644 4140
rect 339552 4100 351644 4128
rect 339552 4088 339558 4100
rect 351638 4088 351644 4100
rect 351696 4088 351702 4140
rect 356054 4088 356060 4140
rect 356112 4128 356118 4140
rect 369394 4128 369400 4140
rect 356112 4100 369400 4128
rect 356112 4088 356118 4100
rect 369394 4088 369400 4100
rect 369452 4088 369458 4140
rect 380986 4088 380992 4140
rect 381044 4128 381050 4140
rect 396534 4128 396540 4140
rect 381044 4100 396540 4128
rect 381044 4088 381050 4100
rect 396534 4088 396540 4100
rect 396592 4088 396598 4140
rect 398834 4088 398840 4140
rect 398892 4128 398898 4140
rect 399110 4128 399116 4140
rect 398892 4100 399116 4128
rect 398892 4088 398898 4100
rect 399110 4088 399116 4100
rect 399168 4088 399174 4140
rect 401686 4088 401692 4140
rect 401744 4128 401750 4140
rect 418982 4128 418988 4140
rect 401744 4100 418988 4128
rect 401744 4088 401750 4100
rect 418982 4088 418988 4100
rect 419040 4088 419046 4140
rect 447134 4088 447140 4140
rect 447192 4128 447198 4140
rect 467466 4128 467472 4140
rect 447192 4100 467472 4128
rect 447192 4088 447198 4100
rect 467466 4088 467472 4100
rect 467524 4088 467530 4140
rect 485038 4088 485044 4140
rect 485096 4128 485102 4140
rect 500586 4128 500592 4140
rect 485096 4100 500592 4128
rect 485096 4088 485102 4100
rect 500586 4088 500592 4100
rect 500644 4088 500650 4140
rect 523126 4088 523132 4140
rect 523184 4128 523190 4140
rect 524322 4128 524328 4140
rect 523184 4100 524328 4128
rect 523184 4088 523190 4100
rect 524322 4088 524328 4100
rect 524380 4088 524386 4140
rect 555418 4088 555424 4140
rect 555476 4128 555482 4140
rect 564434 4128 564440 4140
rect 555476 4100 564440 4128
rect 555476 4088 555482 4100
rect 564434 4088 564440 4100
rect 564492 4088 564498 4140
rect 226426 4020 226432 4072
rect 226484 4060 226490 4072
rect 229830 4060 229836 4072
rect 226484 4032 229836 4060
rect 226484 4020 226490 4032
rect 229830 4020 229836 4032
rect 229888 4020 229894 4072
rect 234706 4020 234712 4072
rect 234764 4060 234770 4072
rect 239306 4060 239312 4072
rect 234764 4032 239312 4060
rect 234764 4020 234770 4032
rect 239306 4020 239312 4032
rect 239364 4020 239370 4072
rect 271966 4020 271972 4072
rect 272024 4060 272030 4072
rect 279510 4060 279516 4072
rect 272024 4032 279516 4060
rect 272024 4020 272030 4032
rect 279510 4020 279516 4032
rect 279568 4020 279574 4072
rect 295334 4020 295340 4072
rect 295392 4060 295398 4072
rect 304350 4060 304356 4072
rect 295392 4032 304356 4060
rect 295392 4020 295398 4032
rect 304350 4020 304356 4032
rect 304408 4020 304414 4072
rect 309778 4020 309784 4072
rect 309836 4060 309842 4072
rect 317322 4060 317328 4072
rect 309836 4032 317328 4060
rect 309836 4020 309842 4032
rect 317322 4020 317328 4032
rect 317380 4020 317386 4072
rect 322934 4020 322940 4072
rect 322992 4060 322998 4072
rect 333882 4060 333888 4072
rect 322992 4032 333888 4060
rect 322992 4020 322998 4032
rect 333882 4020 333888 4032
rect 333940 4020 333946 4072
rect 333974 4020 333980 4072
rect 334032 4060 334038 4072
rect 345750 4060 345756 4072
rect 334032 4032 345756 4060
rect 334032 4020 334038 4032
rect 345750 4020 345756 4032
rect 345808 4020 345814 4072
rect 347774 4020 347780 4072
rect 347832 4060 347838 4072
rect 361114 4060 361120 4072
rect 347832 4032 361120 4060
rect 347832 4020 347838 4032
rect 361114 4020 361120 4032
rect 361172 4020 361178 4072
rect 362954 4020 362960 4072
rect 363012 4060 363018 4072
rect 377674 4060 377680 4072
rect 363012 4032 377680 4060
rect 363012 4020 363018 4032
rect 377674 4020 377680 4032
rect 377732 4020 377738 4072
rect 387886 4020 387892 4072
rect 387944 4060 387950 4072
rect 387944 4032 389174 4060
rect 387944 4020 387950 4032
rect 263594 3952 263600 4004
rect 263652 3992 263658 4004
rect 270034 3992 270040 4004
rect 263652 3964 270040 3992
rect 263652 3952 263658 3964
rect 270034 3952 270040 3964
rect 270092 3952 270098 4004
rect 298094 3952 298100 4004
rect 298152 3992 298158 4004
rect 306742 3992 306748 4004
rect 298152 3964 306748 3992
rect 298152 3952 298158 3964
rect 306742 3952 306748 3964
rect 306800 3952 306806 4004
rect 310514 3952 310520 4004
rect 310572 3992 310578 4004
rect 320910 3992 320916 4004
rect 310572 3964 320916 3992
rect 310572 3952 310578 3964
rect 320910 3952 320916 3964
rect 320968 3952 320974 4004
rect 323578 3952 323584 4004
rect 323636 3992 323642 4004
rect 330386 3992 330392 4004
rect 323636 3964 330392 3992
rect 323636 3952 323642 3964
rect 330386 3952 330392 3964
rect 330444 3952 330450 4004
rect 338114 3952 338120 4004
rect 338172 3992 338178 4004
rect 350442 3992 350448 4004
rect 338172 3964 350448 3992
rect 338172 3952 338178 3964
rect 350442 3952 350448 3964
rect 350500 3952 350506 4004
rect 356238 3952 356244 4004
rect 356296 3992 356302 4004
rect 370590 3992 370596 4004
rect 356296 3964 370596 3992
rect 356296 3952 356302 3964
rect 370590 3952 370596 3964
rect 370648 3952 370654 4004
rect 371234 3952 371240 4004
rect 371292 3992 371298 4004
rect 385954 3992 385960 4004
rect 371292 3964 385960 3992
rect 371292 3952 371298 3964
rect 385954 3952 385960 3964
rect 386012 3952 386018 4004
rect 389146 3992 389174 4032
rect 391934 4020 391940 4072
rect 391992 4060 391998 4072
rect 408402 4060 408408 4072
rect 391992 4032 408408 4060
rect 391992 4020 391998 4032
rect 408402 4020 408408 4032
rect 408460 4020 408466 4072
rect 408586 4020 408592 4072
rect 408644 4060 408650 4072
rect 426158 4060 426164 4072
rect 408644 4032 426164 4060
rect 408644 4020 408650 4032
rect 426158 4020 426164 4032
rect 426216 4020 426222 4072
rect 441614 4020 441620 4072
rect 441672 4060 441678 4072
rect 456058 4060 456064 4072
rect 441672 4032 456064 4060
rect 441672 4020 441678 4032
rect 456058 4020 456064 4032
rect 456116 4020 456122 4072
rect 490558 4020 490564 4072
rect 490616 4060 490622 4072
rect 511258 4060 511264 4072
rect 490616 4032 511264 4060
rect 490616 4020 490622 4032
rect 511258 4020 511264 4032
rect 511316 4020 511322 4072
rect 529198 4020 529204 4072
rect 529256 4060 529262 4072
rect 549070 4060 549076 4072
rect 529256 4032 549076 4060
rect 529256 4020 529262 4032
rect 549070 4020 549076 4032
rect 549128 4020 549134 4072
rect 556798 4020 556804 4072
rect 556856 4060 556862 4072
rect 571518 4060 571524 4072
rect 556856 4032 571524 4060
rect 556856 4020 556862 4032
rect 571518 4020 571524 4032
rect 571576 4020 571582 4072
rect 403618 3992 403624 4004
rect 389146 3964 398834 3992
rect 264238 3884 264244 3936
rect 264296 3924 264302 3936
rect 267734 3924 267740 3936
rect 264296 3896 267740 3924
rect 264296 3884 264302 3896
rect 267734 3884 267740 3896
rect 267792 3884 267798 3936
rect 277486 3884 277492 3936
rect 277544 3924 277550 3936
rect 285398 3924 285404 3936
rect 277544 3896 285404 3924
rect 277544 3884 277550 3896
rect 285398 3884 285404 3896
rect 285456 3884 285462 3936
rect 285674 3884 285680 3936
rect 285732 3924 285738 3936
rect 293678 3924 293684 3936
rect 285732 3896 293684 3924
rect 285732 3884 285738 3896
rect 293678 3884 293684 3896
rect 293736 3884 293742 3936
rect 303614 3884 303620 3936
rect 303672 3924 303678 3936
rect 312630 3924 312636 3936
rect 303672 3896 312636 3924
rect 303672 3884 303678 3896
rect 312630 3884 312636 3896
rect 312688 3884 312694 3936
rect 318794 3884 318800 3936
rect 318852 3924 318858 3936
rect 329190 3924 329196 3936
rect 318852 3896 329196 3924
rect 318852 3884 318858 3896
rect 329190 3884 329196 3896
rect 329248 3884 329254 3936
rect 332594 3884 332600 3936
rect 332652 3924 332658 3936
rect 344554 3924 344560 3936
rect 332652 3896 344560 3924
rect 332652 3884 332658 3896
rect 344554 3884 344560 3896
rect 344612 3884 344618 3936
rect 345014 3884 345020 3936
rect 345072 3924 345078 3936
rect 357526 3924 357532 3936
rect 345072 3896 357532 3924
rect 345072 3884 345078 3896
rect 357526 3884 357532 3896
rect 357584 3884 357590 3936
rect 360194 3884 360200 3936
rect 360252 3924 360258 3936
rect 374086 3924 374092 3936
rect 360252 3896 374092 3924
rect 360252 3884 360258 3896
rect 374086 3884 374092 3896
rect 374144 3884 374150 3936
rect 383746 3884 383752 3936
rect 383804 3924 383810 3936
rect 398806 3924 398834 3964
rect 398944 3964 403624 3992
rect 398944 3924 398972 3964
rect 403618 3952 403624 3964
rect 403676 3952 403682 4004
rect 409966 3952 409972 4004
rect 410024 3992 410030 4004
rect 428458 3992 428464 4004
rect 410024 3964 428464 3992
rect 410024 3952 410030 3964
rect 428458 3952 428464 3964
rect 428516 3952 428522 4004
rect 430758 3952 430764 4004
rect 430816 3992 430822 4004
rect 450906 3992 450912 4004
rect 430816 3964 450912 3992
rect 430816 3952 430822 3964
rect 450906 3952 450912 3964
rect 450964 3952 450970 4004
rect 456978 3952 456984 4004
rect 457036 3992 457042 4004
rect 478138 3992 478144 4004
rect 457036 3964 478144 3992
rect 457036 3952 457042 3964
rect 478138 3952 478144 3964
rect 478196 3952 478202 4004
rect 492674 3952 492680 4004
rect 492732 3992 492738 4004
rect 517146 3992 517152 4004
rect 492732 3964 517152 3992
rect 492732 3952 492738 3964
rect 517146 3952 517152 3964
rect 517204 3952 517210 4004
rect 522298 3952 522304 4004
rect 522356 3992 522362 4004
rect 545482 3992 545488 4004
rect 522356 3964 545488 3992
rect 522356 3952 522362 3964
rect 545482 3952 545488 3964
rect 545540 3952 545546 4004
rect 560938 3952 560944 4004
rect 560996 3992 561002 4004
rect 582190 3992 582196 4004
rect 560996 3964 582196 3992
rect 560996 3952 561002 3964
rect 582190 3952 582196 3964
rect 582248 3952 582254 4004
rect 383804 3896 389174 3924
rect 398806 3896 398972 3924
rect 383804 3884 383810 3896
rect 102226 3816 102232 3868
rect 102284 3856 102290 3868
rect 105538 3856 105544 3868
rect 102284 3828 105544 3856
rect 102284 3816 102290 3828
rect 105538 3816 105544 3828
rect 105596 3816 105602 3868
rect 227806 3816 227812 3868
rect 227864 3856 227870 3868
rect 231026 3856 231032 3868
rect 227864 3828 231032 3856
rect 227864 3816 227870 3828
rect 231026 3816 231032 3828
rect 231084 3816 231090 3868
rect 247034 3816 247040 3868
rect 247092 3856 247098 3868
rect 252370 3856 252376 3868
rect 247092 3828 252376 3856
rect 247092 3816 247098 3828
rect 252370 3816 252376 3828
rect 252428 3816 252434 3868
rect 281626 3816 281632 3868
rect 281684 3856 281690 3868
rect 290182 3856 290188 3868
rect 281684 3828 290188 3856
rect 281684 3816 281690 3828
rect 290182 3816 290188 3828
rect 290240 3816 290246 3868
rect 306374 3816 306380 3868
rect 306432 3856 306438 3868
rect 316218 3856 316224 3868
rect 306432 3828 316224 3856
rect 306432 3816 306438 3828
rect 316218 3816 316224 3828
rect 316276 3816 316282 3868
rect 317414 3816 317420 3868
rect 317472 3856 317478 3868
rect 327994 3856 328000 3868
rect 317472 3828 328000 3856
rect 317472 3816 317478 3828
rect 327994 3816 328000 3828
rect 328052 3816 328058 3868
rect 329834 3816 329840 3868
rect 329892 3856 329898 3868
rect 342162 3856 342168 3868
rect 329892 3828 342168 3856
rect 329892 3816 329898 3828
rect 342162 3816 342168 3828
rect 342220 3816 342226 3868
rect 354674 3816 354680 3868
rect 354732 3856 354738 3868
rect 368198 3856 368204 3868
rect 354732 3828 368204 3856
rect 354732 3816 354738 3828
rect 368198 3816 368204 3828
rect 368256 3816 368262 3868
rect 368474 3816 368480 3868
rect 368532 3856 368538 3868
rect 383562 3856 383568 3868
rect 368532 3828 383568 3856
rect 368532 3816 368538 3828
rect 383562 3816 383568 3828
rect 383620 3816 383626 3868
rect 389146 3856 389174 3896
rect 399110 3884 399116 3936
rect 399168 3924 399174 3936
rect 415486 3924 415492 3936
rect 399168 3896 415492 3924
rect 399168 3884 399174 3896
rect 415486 3884 415492 3896
rect 415544 3884 415550 3936
rect 423674 3884 423680 3936
rect 423732 3924 423738 3936
rect 442626 3924 442632 3936
rect 423732 3896 442632 3924
rect 423732 3884 423738 3896
rect 442626 3884 442632 3896
rect 442684 3884 442690 3936
rect 447226 3884 447232 3936
rect 447284 3924 447290 3936
rect 468662 3924 468668 3936
rect 447284 3896 468668 3924
rect 447284 3884 447290 3896
rect 468662 3884 468668 3896
rect 468720 3884 468726 3936
rect 486418 3884 486424 3936
rect 486476 3924 486482 3936
rect 504174 3924 504180 3936
rect 486476 3896 504180 3924
rect 486476 3884 486482 3896
rect 504174 3884 504180 3896
rect 504232 3884 504238 3936
rect 506566 3884 506572 3936
rect 506624 3924 506630 3936
rect 532510 3924 532516 3936
rect 506624 3896 532516 3924
rect 506624 3884 506630 3896
rect 532510 3884 532516 3896
rect 532568 3884 532574 3936
rect 556890 3884 556896 3936
rect 556948 3924 556954 3936
rect 578602 3924 578608 3936
rect 556948 3896 578608 3924
rect 556948 3884 556954 3896
rect 578602 3884 578608 3896
rect 578660 3884 578666 3936
rect 400122 3856 400128 3868
rect 389146 3828 400128 3856
rect 400122 3816 400128 3828
rect 400180 3816 400186 3868
rect 416774 3816 416780 3868
rect 416832 3856 416838 3868
rect 435542 3856 435548 3868
rect 416832 3828 435548 3856
rect 416832 3816 416838 3828
rect 435542 3816 435548 3828
rect 435600 3816 435606 3868
rect 452654 3816 452660 3868
rect 452712 3856 452718 3868
rect 474550 3856 474556 3868
rect 452712 3828 474556 3856
rect 452712 3816 452718 3828
rect 474550 3816 474556 3828
rect 474608 3816 474614 3868
rect 499574 3816 499580 3868
rect 499632 3856 499638 3868
rect 524230 3856 524236 3868
rect 499632 3828 524236 3856
rect 499632 3816 499638 3828
rect 524230 3816 524236 3828
rect 524288 3816 524294 3868
rect 524322 3816 524328 3868
rect 524380 3856 524386 3868
rect 550266 3856 550272 3868
rect 524380 3828 550272 3856
rect 524380 3816 524386 3828
rect 550266 3816 550272 3828
rect 550324 3816 550330 3868
rect 551278 3816 551284 3868
rect 551336 3856 551342 3868
rect 577406 3856 577412 3868
rect 551336 3828 577412 3856
rect 551336 3816 551342 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 121086 3748 121092 3800
rect 121144 3788 121150 3800
rect 124858 3788 124864 3800
rect 121144 3760 124864 3788
rect 121144 3748 121150 3760
rect 124858 3748 124864 3760
rect 124916 3748 124922 3800
rect 256694 3748 256700 3800
rect 256752 3788 256758 3800
rect 262950 3788 262956 3800
rect 256752 3760 262956 3788
rect 256752 3748 256758 3760
rect 262950 3748 262956 3760
rect 263008 3748 263014 3800
rect 282914 3748 282920 3800
rect 282972 3788 282978 3800
rect 291378 3788 291384 3800
rect 282972 3760 291384 3788
rect 282972 3748 282978 3760
rect 291378 3748 291384 3760
rect 291436 3748 291442 3800
rect 299474 3748 299480 3800
rect 299532 3788 299538 3800
rect 309042 3788 309048 3800
rect 299532 3760 309048 3788
rect 299532 3748 299538 3760
rect 309042 3748 309048 3760
rect 309100 3748 309106 3800
rect 311894 3748 311900 3800
rect 311952 3788 311958 3800
rect 322106 3788 322112 3800
rect 311952 3760 322112 3788
rect 311952 3748 311958 3760
rect 322106 3748 322112 3760
rect 322164 3748 322170 3800
rect 328454 3748 328460 3800
rect 328512 3788 328518 3800
rect 339862 3788 339868 3800
rect 328512 3760 339868 3788
rect 328512 3748 328518 3760
rect 339862 3748 339868 3760
rect 339920 3748 339926 3800
rect 343634 3748 343640 3800
rect 343692 3788 343698 3800
rect 356330 3788 356336 3800
rect 343692 3760 356336 3788
rect 343692 3748 343698 3760
rect 356330 3748 356336 3760
rect 356388 3748 356394 3800
rect 357434 3748 357440 3800
rect 357492 3788 357498 3800
rect 357492 3760 362448 3788
rect 357492 3748 357498 3760
rect 6886 3692 16574 3720
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 6886 3584 6914 3692
rect 2924 3556 6914 3584
rect 2924 3544 2930 3556
rect 15286 3544 15292 3596
rect 15344 3544 15350 3596
rect 16546 3584 16574 3692
rect 237466 3680 237472 3732
rect 237524 3720 237530 3732
rect 241698 3720 241704 3732
rect 237524 3692 241704 3720
rect 237524 3680 237530 3692
rect 241698 3680 241704 3692
rect 241756 3680 241762 3732
rect 249978 3680 249984 3732
rect 250036 3720 250042 3732
rect 255866 3720 255872 3732
rect 250036 3692 255872 3720
rect 250036 3680 250042 3692
rect 255866 3680 255872 3692
rect 255924 3680 255930 3732
rect 266354 3680 266360 3732
rect 266412 3720 266418 3732
rect 272426 3720 272432 3732
rect 266412 3692 272432 3720
rect 266412 3680 266418 3692
rect 272426 3680 272432 3692
rect 272484 3680 272490 3732
rect 273254 3680 273260 3732
rect 273312 3720 273318 3732
rect 280706 3720 280712 3732
rect 273312 3692 280712 3720
rect 273312 3680 273318 3692
rect 280706 3680 280712 3692
rect 280764 3680 280770 3732
rect 304994 3680 305000 3732
rect 305052 3720 305058 3732
rect 315022 3720 315028 3732
rect 305052 3692 315028 3720
rect 305052 3680 305058 3692
rect 315022 3680 315028 3692
rect 315080 3680 315086 3732
rect 316034 3680 316040 3732
rect 316092 3720 316098 3732
rect 326798 3720 326804 3732
rect 316092 3692 326804 3720
rect 316092 3680 316098 3692
rect 326798 3680 326804 3692
rect 326856 3680 326862 3732
rect 327074 3680 327080 3732
rect 327132 3720 327138 3732
rect 338666 3720 338672 3732
rect 327132 3692 338672 3720
rect 327132 3680 327138 3692
rect 338666 3680 338672 3692
rect 338724 3680 338730 3732
rect 349154 3680 349160 3732
rect 349212 3720 349218 3732
rect 362310 3720 362316 3732
rect 349212 3692 362316 3720
rect 349212 3680 349218 3692
rect 362310 3680 362316 3692
rect 362368 3680 362374 3732
rect 362420 3720 362448 3760
rect 364334 3748 364340 3800
rect 364392 3788 364398 3800
rect 378870 3788 378876 3800
rect 364392 3760 378876 3788
rect 364392 3748 364398 3760
rect 378870 3748 378876 3760
rect 378928 3748 378934 3800
rect 397454 3748 397460 3800
rect 397512 3788 397518 3800
rect 414290 3788 414296 3800
rect 397512 3760 414296 3788
rect 397512 3748 397518 3760
rect 414290 3748 414296 3760
rect 414348 3748 414354 3800
rect 418154 3748 418160 3800
rect 418212 3788 418218 3800
rect 436738 3788 436744 3800
rect 418212 3760 436744 3788
rect 418212 3748 418218 3760
rect 436738 3748 436744 3760
rect 436796 3748 436802 3800
rect 439498 3748 439504 3800
rect 439556 3788 439562 3800
rect 446214 3788 446220 3800
rect 439556 3760 446220 3788
rect 439556 3748 439562 3760
rect 446214 3748 446220 3760
rect 446272 3748 446278 3800
rect 449894 3748 449900 3800
rect 449952 3788 449958 3800
rect 471054 3788 471060 3800
rect 449952 3760 471060 3788
rect 449952 3748 449958 3760
rect 471054 3748 471060 3760
rect 471112 3748 471118 3800
rect 482278 3748 482284 3800
rect 482336 3788 482342 3800
rect 497090 3788 497096 3800
rect 482336 3760 497096 3788
rect 482336 3748 482342 3760
rect 497090 3748 497096 3760
rect 497148 3748 497154 3800
rect 499758 3748 499764 3800
rect 499816 3788 499822 3800
rect 525426 3788 525432 3800
rect 499816 3760 525432 3788
rect 499816 3748 499822 3760
rect 525426 3748 525432 3760
rect 525484 3748 525490 3800
rect 525886 3748 525892 3800
rect 525944 3788 525950 3800
rect 553762 3788 553768 3800
rect 525944 3760 553768 3788
rect 525944 3748 525950 3760
rect 553762 3748 553768 3760
rect 553820 3748 553826 3800
rect 558178 3748 558184 3800
rect 558236 3788 558242 3800
rect 580994 3788 581000 3800
rect 558236 3760 581000 3788
rect 558236 3748 558242 3760
rect 580994 3748 581000 3760
rect 581052 3748 581058 3800
rect 362420 3692 367140 3720
rect 209774 3612 209780 3664
rect 209832 3652 209838 3664
rect 212166 3652 212172 3664
rect 209832 3624 212172 3652
rect 209832 3612 209838 3624
rect 212166 3612 212172 3624
rect 212224 3612 212230 3664
rect 212626 3612 212632 3664
rect 212684 3652 212690 3664
rect 215662 3652 215668 3664
rect 212684 3624 215668 3652
rect 212684 3612 212690 3624
rect 215662 3612 215668 3624
rect 215720 3612 215726 3664
rect 276014 3612 276020 3664
rect 276072 3652 276078 3664
rect 283098 3652 283104 3664
rect 276072 3624 283104 3652
rect 276072 3612 276078 3624
rect 283098 3612 283104 3624
rect 283156 3612 283162 3664
rect 284294 3612 284300 3664
rect 284352 3652 284358 3664
rect 292574 3652 292580 3664
rect 284352 3624 292580 3652
rect 284352 3612 284358 3624
rect 292574 3612 292580 3624
rect 292632 3612 292638 3664
rect 293954 3612 293960 3664
rect 294012 3652 294018 3664
rect 303154 3652 303160 3664
rect 294012 3624 303160 3652
rect 294012 3612 294018 3624
rect 303154 3612 303160 3624
rect 303212 3612 303218 3664
rect 307754 3612 307760 3664
rect 307812 3652 307818 3664
rect 318518 3652 318524 3664
rect 307812 3624 318524 3652
rect 307812 3612 307818 3624
rect 318518 3612 318524 3624
rect 318576 3612 318582 3664
rect 320174 3612 320180 3664
rect 320232 3652 320238 3664
rect 331582 3652 331588 3664
rect 320232 3624 331588 3652
rect 320232 3612 320238 3624
rect 331582 3612 331588 3624
rect 331640 3612 331646 3664
rect 335354 3612 335360 3664
rect 335412 3652 335418 3664
rect 346946 3652 346952 3664
rect 335412 3624 346952 3652
rect 335412 3612 335418 3624
rect 346946 3612 346952 3624
rect 347004 3612 347010 3664
rect 351914 3612 351920 3664
rect 351972 3652 351978 3664
rect 365806 3652 365812 3664
rect 351972 3624 365812 3652
rect 351972 3612 351978 3624
rect 365806 3612 365812 3624
rect 365864 3612 365870 3664
rect 367112 3652 367140 3692
rect 367186 3680 367192 3732
rect 367244 3720 367250 3732
rect 382366 3720 382372 3732
rect 367244 3692 382372 3720
rect 367244 3680 367250 3692
rect 382366 3680 382372 3692
rect 382424 3680 382430 3732
rect 385034 3680 385040 3732
rect 385092 3720 385098 3732
rect 401318 3720 401324 3732
rect 385092 3692 401324 3720
rect 385092 3680 385098 3692
rect 401318 3680 401324 3692
rect 401376 3680 401382 3732
rect 411898 3720 411904 3732
rect 403636 3692 411904 3720
rect 371694 3652 371700 3664
rect 367112 3624 371700 3652
rect 371694 3612 371700 3624
rect 371752 3612 371758 3664
rect 375466 3612 375472 3664
rect 375524 3652 375530 3664
rect 390554 3652 390560 3664
rect 375524 3624 390560 3652
rect 375524 3612 375530 3624
rect 390554 3612 390560 3624
rect 390612 3612 390618 3664
rect 390646 3612 390652 3664
rect 390704 3652 390710 3664
rect 402974 3652 402980 3664
rect 390704 3624 402980 3652
rect 390704 3612 390710 3624
rect 402974 3612 402980 3624
rect 403032 3612 403038 3664
rect 16666 3584 16672 3596
rect 16546 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 130562 3544 130568 3596
rect 130620 3584 130626 3596
rect 133966 3584 133972 3596
rect 130620 3556 133972 3584
rect 130620 3544 130626 3556
rect 133966 3544 133972 3556
rect 134024 3544 134030 3596
rect 138842 3544 138848 3596
rect 138900 3584 138906 3596
rect 142246 3584 142252 3596
rect 138900 3556 142252 3584
rect 138900 3544 138906 3556
rect 142246 3544 142252 3556
rect 142304 3544 142310 3596
rect 143626 3544 143632 3596
rect 143684 3584 143690 3596
rect 144730 3584 144736 3596
rect 143684 3556 144736 3584
rect 143684 3544 143690 3556
rect 144730 3544 144736 3556
rect 144788 3544 144794 3596
rect 191926 3544 191932 3596
rect 191984 3584 191990 3596
rect 193214 3584 193220 3596
rect 191984 3556 193220 3584
rect 191984 3544 191990 3556
rect 193214 3544 193220 3556
rect 193272 3544 193278 3596
rect 197446 3544 197452 3596
rect 197504 3584 197510 3596
rect 199102 3584 199108 3596
rect 197504 3556 199108 3584
rect 197504 3544 197510 3556
rect 199102 3544 199108 3556
rect 199160 3544 199166 3596
rect 200206 3544 200212 3596
rect 200264 3584 200270 3596
rect 201494 3584 201500 3596
rect 200264 3556 201500 3584
rect 200264 3544 200270 3556
rect 201494 3544 201500 3556
rect 201552 3544 201558 3596
rect 204346 3544 204352 3596
rect 204404 3584 204410 3596
rect 206186 3584 206192 3596
rect 204404 3556 206192 3584
rect 204404 3544 204410 3556
rect 206186 3544 206192 3556
rect 206244 3544 206250 3596
rect 207014 3544 207020 3596
rect 207072 3584 207078 3596
rect 207072 3556 209774 3584
rect 207072 3544 207078 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 15304 3516 15332 3544
rect 209746 3528 209774 3556
rect 214006 3544 214012 3596
rect 214064 3584 214070 3596
rect 216858 3584 216864 3596
rect 214064 3556 216864 3584
rect 214064 3544 214070 3556
rect 216858 3544 216864 3556
rect 216916 3544 216922 3596
rect 218054 3544 218060 3596
rect 218112 3584 218118 3596
rect 220446 3584 220452 3596
rect 218112 3556 220452 3584
rect 218112 3544 218118 3556
rect 220446 3544 220452 3556
rect 220504 3544 220510 3596
rect 223574 3544 223580 3596
rect 223632 3584 223638 3596
rect 227530 3584 227536 3596
rect 223632 3556 227536 3584
rect 223632 3544 223638 3556
rect 227530 3544 227536 3556
rect 227588 3544 227594 3596
rect 233326 3544 233332 3596
rect 233384 3584 233390 3596
rect 237006 3584 237012 3596
rect 233384 3556 237012 3584
rect 233384 3544 233390 3556
rect 237006 3544 237012 3556
rect 237064 3544 237070 3596
rect 244274 3544 244280 3596
rect 244332 3584 244338 3596
rect 249978 3584 249984 3596
rect 244332 3556 249984 3584
rect 244332 3544 244338 3556
rect 249978 3544 249984 3556
rect 250036 3544 250042 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 257062 3584 257068 3596
rect 251232 3556 257068 3584
rect 251232 3544 251238 3556
rect 257062 3544 257068 3556
rect 257120 3544 257126 3596
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 265342 3584 265348 3596
rect 259512 3556 265348 3584
rect 259512 3544 259518 3556
rect 265342 3544 265348 3556
rect 265400 3544 265406 3596
rect 266446 3544 266452 3596
rect 266504 3584 266510 3596
rect 273622 3584 273628 3596
rect 266504 3556 273628 3584
rect 266504 3544 266510 3556
rect 273622 3544 273628 3556
rect 273680 3544 273686 3596
rect 274634 3544 274640 3596
rect 274692 3584 274698 3596
rect 281902 3584 281908 3596
rect 274692 3556 281908 3584
rect 274692 3544 274698 3556
rect 281902 3544 281908 3556
rect 281960 3544 281966 3596
rect 287146 3544 287152 3596
rect 287204 3584 287210 3596
rect 294874 3584 294880 3596
rect 287204 3556 294880 3584
rect 287204 3544 287210 3556
rect 294874 3544 294880 3556
rect 294932 3544 294938 3596
rect 303706 3544 303712 3596
rect 303764 3584 303770 3596
rect 313826 3584 313832 3596
rect 303764 3556 313832 3584
rect 303764 3544 303770 3556
rect 313826 3544 313832 3556
rect 313884 3544 313890 3596
rect 314654 3544 314660 3596
rect 314712 3584 314718 3596
rect 325602 3584 325608 3596
rect 314712 3556 325608 3584
rect 314712 3544 314718 3556
rect 325602 3544 325608 3556
rect 325660 3544 325666 3596
rect 325694 3544 325700 3596
rect 325752 3584 325758 3596
rect 337470 3584 337476 3596
rect 325752 3556 337476 3584
rect 325752 3544 325758 3556
rect 337470 3544 337476 3556
rect 337528 3544 337534 3596
rect 342254 3544 342260 3596
rect 342312 3584 342318 3596
rect 355226 3584 355232 3596
rect 342312 3556 355232 3584
rect 342312 3544 342318 3556
rect 355226 3544 355232 3556
rect 355284 3544 355290 3596
rect 358814 3544 358820 3596
rect 358872 3584 358878 3596
rect 372890 3584 372896 3596
rect 358872 3556 372896 3584
rect 358872 3544 358878 3556
rect 372890 3544 372896 3556
rect 372948 3544 372954 3596
rect 373994 3544 374000 3596
rect 374052 3584 374058 3596
rect 389450 3584 389456 3596
rect 374052 3556 389456 3584
rect 374052 3544 374058 3556
rect 389450 3544 389456 3556
rect 389508 3544 389514 3596
rect 394786 3544 394792 3596
rect 394844 3584 394850 3596
rect 403636 3584 403664 3692
rect 411898 3680 411904 3692
rect 411956 3680 411962 3732
rect 421374 3720 421380 3732
rect 412606 3692 421380 3720
rect 404354 3612 404360 3664
rect 404412 3652 404418 3664
rect 412606 3652 412634 3692
rect 421374 3680 421380 3692
rect 421432 3680 421438 3732
rect 425054 3680 425060 3732
rect 425112 3720 425118 3732
rect 443822 3720 443828 3732
rect 425112 3692 443828 3720
rect 425112 3680 425118 3692
rect 443822 3680 443828 3692
rect 443880 3680 443886 3732
rect 456058 3680 456064 3732
rect 456116 3720 456122 3732
rect 461578 3720 461584 3732
rect 456116 3692 461584 3720
rect 456116 3680 456122 3692
rect 461578 3680 461584 3692
rect 461636 3680 461642 3732
rect 463694 3680 463700 3732
rect 463752 3720 463758 3732
rect 486418 3720 486424 3732
rect 463752 3692 486424 3720
rect 463752 3680 463758 3692
rect 486418 3680 486424 3692
rect 486476 3680 486482 3732
rect 503714 3680 503720 3732
rect 503772 3720 503778 3732
rect 529014 3720 529020 3732
rect 503772 3692 529020 3720
rect 503772 3680 503778 3692
rect 529014 3680 529020 3692
rect 529072 3680 529078 3732
rect 532786 3680 532792 3732
rect 532844 3720 532850 3732
rect 560846 3720 560852 3732
rect 532844 3692 560852 3720
rect 532844 3680 532850 3692
rect 560846 3680 560852 3692
rect 560904 3680 560910 3732
rect 566458 3680 566464 3732
rect 566516 3720 566522 3732
rect 576302 3720 576308 3732
rect 566516 3692 576308 3720
rect 566516 3680 566522 3692
rect 576302 3680 576308 3692
rect 576360 3680 576366 3732
rect 404412 3624 412634 3652
rect 404412 3612 404418 3624
rect 414014 3612 414020 3664
rect 414072 3652 414078 3664
rect 433242 3652 433248 3664
rect 414072 3624 433248 3652
rect 414072 3612 414078 3624
rect 433242 3612 433248 3624
rect 433300 3612 433306 3664
rect 434714 3612 434720 3664
rect 434772 3652 434778 3664
rect 454494 3652 454500 3664
rect 434772 3624 454500 3652
rect 434772 3612 434778 3624
rect 454494 3612 454500 3624
rect 454552 3612 454558 3664
rect 456794 3612 456800 3664
rect 456852 3652 456858 3664
rect 458266 3652 458272 3664
rect 456852 3624 458272 3652
rect 456852 3612 456858 3624
rect 458266 3612 458272 3624
rect 458324 3612 458330 3664
rect 460934 3612 460940 3664
rect 460992 3652 460998 3664
rect 482830 3652 482836 3664
rect 460992 3624 482836 3652
rect 460992 3612 460998 3624
rect 482830 3612 482836 3624
rect 482888 3612 482894 3664
rect 483106 3612 483112 3664
rect 483164 3652 483170 3664
rect 507670 3652 507676 3664
rect 483164 3624 507676 3652
rect 483164 3612 483170 3624
rect 507670 3612 507676 3624
rect 507728 3612 507734 3664
rect 510614 3612 510620 3664
rect 510672 3652 510678 3664
rect 536098 3652 536104 3664
rect 510672 3624 536104 3652
rect 510672 3612 510678 3624
rect 536098 3612 536104 3624
rect 536156 3612 536162 3664
rect 539686 3612 539692 3664
rect 539744 3652 539750 3664
rect 568022 3652 568028 3664
rect 539744 3624 568028 3652
rect 539744 3612 539750 3624
rect 568022 3612 568028 3624
rect 568080 3612 568086 3664
rect 410794 3584 410800 3596
rect 394844 3556 403664 3584
rect 405016 3556 410800 3584
rect 394844 3544 394850 3556
rect 1728 3488 15332 3516
rect 1728 3476 1734 3488
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 28534 3516 28540 3528
rect 27672 3488 28540 3516
rect 27672 3476 27678 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 68278 3516 68284 3528
rect 66772 3488 68284 3516
rect 66772 3476 66778 3488
rect 68278 3476 68284 3488
rect 68336 3476 68342 3528
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 69934 3516 69940 3528
rect 69072 3488 69940 3516
rect 69072 3476 69078 3488
rect 69934 3476 69940 3488
rect 69992 3476 69998 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111610 3516 111616 3528
rect 110564 3488 111616 3516
rect 110564 3476 110570 3488
rect 111610 3476 111616 3488
rect 111668 3476 111674 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119890 3516 119896 3528
rect 118844 3488 119896 3516
rect 118844 3476 118850 3488
rect 119890 3476 119896 3488
rect 119948 3476 119954 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128170 3516 128176 3528
rect 127032 3488 128176 3516
rect 127032 3476 127038 3488
rect 128170 3476 128176 3488
rect 128228 3476 128234 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 169754 3476 169760 3528
rect 169812 3516 169818 3528
rect 170398 3516 170404 3528
rect 169812 3488 170404 3516
rect 169812 3476 169818 3488
rect 170398 3476 170404 3488
rect 170456 3476 170462 3528
rect 172514 3476 172520 3528
rect 172572 3516 172578 3528
rect 172790 3516 172796 3528
rect 172572 3488 172796 3516
rect 172572 3476 172578 3488
rect 172790 3476 172796 3488
rect 172848 3476 172854 3528
rect 179046 3476 179052 3528
rect 179104 3516 179110 3528
rect 179506 3516 179512 3528
rect 179104 3488 179512 3516
rect 179104 3476 179110 3488
rect 179506 3476 179512 3488
rect 179564 3476 179570 3528
rect 186314 3476 186320 3528
rect 186372 3516 186378 3528
rect 186958 3516 186964 3528
rect 186372 3488 186964 3516
rect 186372 3476 186378 3488
rect 186958 3476 186964 3488
rect 187016 3476 187022 3528
rect 205634 3476 205640 3528
rect 205692 3516 205698 3528
rect 207382 3516 207388 3528
rect 205692 3488 207388 3516
rect 205692 3476 205698 3488
rect 207382 3476 207388 3488
rect 207440 3476 207446 3528
rect 209746 3488 209780 3528
rect 209774 3476 209780 3488
rect 209832 3476 209838 3528
rect 216674 3476 216680 3528
rect 216732 3516 216738 3528
rect 219250 3516 219256 3528
rect 216732 3488 219256 3516
rect 216732 3476 216738 3488
rect 219250 3476 219256 3488
rect 219308 3476 219314 3528
rect 220078 3476 220084 3528
rect 220136 3516 220142 3528
rect 221550 3516 221556 3528
rect 220136 3488 221556 3516
rect 220136 3476 220142 3488
rect 221550 3476 221556 3488
rect 221608 3476 221614 3528
rect 222194 3476 222200 3528
rect 222252 3516 222258 3528
rect 225138 3516 225144 3528
rect 222252 3488 225144 3516
rect 222252 3476 222258 3488
rect 225138 3476 225144 3488
rect 225196 3476 225202 3528
rect 231946 3476 231952 3528
rect 232004 3516 232010 3528
rect 235810 3516 235816 3528
rect 232004 3488 235816 3516
rect 232004 3476 232010 3488
rect 235810 3476 235816 3488
rect 235868 3476 235874 3528
rect 240778 3476 240784 3528
rect 240836 3516 240842 3528
rect 244090 3516 244096 3528
rect 240836 3488 244096 3516
rect 240836 3476 240842 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 246298 3476 246304 3528
rect 246356 3516 246362 3528
rect 247586 3516 247592 3528
rect 246356 3488 247592 3516
rect 246356 3476 246362 3488
rect 247586 3476 247592 3488
rect 247644 3476 247650 3528
rect 249794 3476 249800 3528
rect 249852 3516 249858 3528
rect 254670 3516 254676 3528
rect 249852 3488 254676 3516
rect 249852 3476 249858 3488
rect 254670 3476 254676 3488
rect 254728 3476 254734 3528
rect 255314 3476 255320 3528
rect 255372 3516 255378 3528
rect 261754 3516 261760 3528
rect 255372 3488 261760 3516
rect 255372 3476 255378 3488
rect 261754 3476 261760 3488
rect 261812 3476 261818 3528
rect 270586 3476 270592 3528
rect 270644 3516 270650 3528
rect 277118 3516 277124 3528
rect 270644 3488 277124 3516
rect 270644 3476 270650 3488
rect 277118 3476 277124 3488
rect 277176 3476 277182 3528
rect 291194 3476 291200 3528
rect 291252 3516 291258 3528
rect 299658 3516 299664 3528
rect 291252 3488 299664 3516
rect 291252 3476 291258 3488
rect 299658 3476 299664 3488
rect 299716 3476 299722 3528
rect 309134 3476 309140 3528
rect 309192 3516 309198 3528
rect 319714 3516 319720 3528
rect 309192 3488 319720 3516
rect 309192 3476 309198 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 321554 3476 321560 3528
rect 321612 3516 321618 3528
rect 332686 3516 332692 3528
rect 321612 3488 332692 3516
rect 321612 3476 321618 3488
rect 332686 3476 332692 3488
rect 332744 3476 332750 3528
rect 335446 3476 335452 3528
rect 335504 3516 335510 3528
rect 348050 3516 348056 3528
rect 335504 3488 348056 3516
rect 335504 3476 335510 3488
rect 348050 3476 348056 3488
rect 348108 3476 348114 3528
rect 350534 3476 350540 3528
rect 350592 3516 350598 3528
rect 350592 3488 354674 3516
rect 350592 3476 350598 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 13814 3448 13820 3460
rect 624 3420 13820 3448
rect 624 3408 630 3420
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 42886 3448 42892 3460
rect 31352 3420 42892 3448
rect 31352 3408 31358 3420
rect 42886 3408 42892 3420
rect 42944 3408 42950 3460
rect 220814 3408 220820 3460
rect 220872 3448 220878 3460
rect 223942 3448 223948 3460
rect 220872 3420 223948 3448
rect 220872 3408 220878 3420
rect 223942 3408 223948 3420
rect 224000 3408 224006 3460
rect 240226 3408 240232 3460
rect 240284 3448 240290 3460
rect 245194 3448 245200 3460
rect 240284 3420 245200 3448
rect 240284 3408 240290 3420
rect 245194 3408 245200 3420
rect 245252 3408 245258 3460
rect 245654 3408 245660 3460
rect 245712 3448 245718 3460
rect 251174 3448 251180 3460
rect 245712 3420 251180 3448
rect 245712 3408 245718 3420
rect 251174 3408 251180 3420
rect 251232 3408 251238 3460
rect 260834 3408 260840 3460
rect 260892 3448 260898 3460
rect 266538 3448 266544 3460
rect 260892 3420 266544 3448
rect 260892 3408 260898 3420
rect 266538 3408 266544 3420
rect 266596 3408 266602 3460
rect 269114 3408 269120 3460
rect 269172 3448 269178 3460
rect 276014 3448 276020 3460
rect 269172 3420 276020 3448
rect 269172 3408 269178 3420
rect 276014 3408 276020 3420
rect 276072 3408 276078 3460
rect 276106 3408 276112 3460
rect 276164 3448 276170 3460
rect 284294 3448 284300 3460
rect 276164 3420 284300 3448
rect 276164 3408 276170 3420
rect 284294 3408 284300 3420
rect 284352 3408 284358 3460
rect 288434 3408 288440 3460
rect 288492 3448 288498 3460
rect 297266 3448 297272 3460
rect 288492 3420 297272 3448
rect 288492 3408 288498 3420
rect 297266 3408 297272 3420
rect 297324 3408 297330 3460
rect 298186 3408 298192 3460
rect 298244 3448 298250 3460
rect 307938 3448 307944 3460
rect 298244 3420 307944 3448
rect 298244 3408 298250 3420
rect 307938 3408 307944 3420
rect 307996 3408 308002 3460
rect 324498 3408 324504 3460
rect 324556 3448 324562 3460
rect 336274 3448 336280 3460
rect 324556 3420 336280 3448
rect 324556 3408 324562 3420
rect 336274 3408 336280 3420
rect 336332 3408 336338 3460
rect 336734 3408 336740 3460
rect 336792 3448 336798 3460
rect 349246 3448 349252 3460
rect 336792 3420 349252 3448
rect 336792 3408 336798 3420
rect 349246 3408 349252 3420
rect 349304 3408 349310 3460
rect 354646 3448 354674 3488
rect 358078 3476 358084 3528
rect 358136 3516 358142 3528
rect 359918 3516 359924 3528
rect 358136 3488 359924 3516
rect 358136 3476 358142 3488
rect 359918 3476 359924 3488
rect 359976 3476 359982 3528
rect 362218 3476 362224 3528
rect 362276 3516 362282 3528
rect 363506 3516 363512 3528
rect 362276 3488 363512 3516
rect 362276 3476 362282 3488
rect 363506 3476 363512 3488
rect 363564 3476 363570 3528
rect 365714 3476 365720 3528
rect 365772 3516 365778 3528
rect 379974 3516 379980 3528
rect 365772 3488 379980 3516
rect 365772 3476 365778 3488
rect 379974 3476 379980 3488
rect 380032 3476 380038 3528
rect 385678 3476 385684 3528
rect 385736 3516 385742 3528
rect 387150 3516 387156 3528
rect 385736 3488 387156 3516
rect 385736 3476 385742 3488
rect 387150 3476 387156 3488
rect 387208 3476 387214 3528
rect 388070 3476 388076 3528
rect 388128 3516 388134 3528
rect 404814 3516 404820 3528
rect 388128 3488 404820 3516
rect 388128 3476 388134 3488
rect 404814 3476 404820 3488
rect 404872 3476 404878 3528
rect 364610 3448 364616 3460
rect 354646 3420 364616 3448
rect 364610 3408 364616 3420
rect 364668 3408 364674 3460
rect 366358 3408 366364 3460
rect 366416 3448 366422 3460
rect 375282 3448 375288 3460
rect 366416 3420 375288 3448
rect 366416 3408 366422 3420
rect 375282 3408 375288 3420
rect 375340 3408 375346 3460
rect 382274 3408 382280 3460
rect 382332 3448 382338 3460
rect 397730 3448 397736 3460
rect 382332 3420 397736 3448
rect 382332 3408 382338 3420
rect 397730 3408 397736 3420
rect 397788 3408 397794 3460
rect 126974 3340 126980 3392
rect 127032 3380 127038 3392
rect 130470 3380 130476 3392
rect 127032 3352 130476 3380
rect 127032 3340 127038 3352
rect 130470 3340 130476 3352
rect 130528 3340 130534 3392
rect 219434 3340 219440 3392
rect 219492 3380 219498 3392
rect 222746 3380 222752 3392
rect 219492 3352 222752 3380
rect 219492 3340 219498 3352
rect 222746 3340 222752 3352
rect 222804 3340 222810 3392
rect 241514 3340 241520 3392
rect 241572 3380 241578 3392
rect 246390 3380 246396 3392
rect 241572 3352 246396 3380
rect 241572 3340 241578 3352
rect 246390 3340 246396 3352
rect 246448 3340 246454 3392
rect 248414 3340 248420 3392
rect 248472 3380 248478 3392
rect 253474 3380 253480 3392
rect 248472 3352 253480 3380
rect 248472 3340 248478 3352
rect 253474 3340 253480 3352
rect 253532 3340 253538 3392
rect 258074 3340 258080 3392
rect 258132 3380 258138 3392
rect 264146 3380 264152 3392
rect 258132 3352 264152 3380
rect 258132 3340 258138 3352
rect 264146 3340 264152 3352
rect 264204 3340 264210 3392
rect 267826 3340 267832 3392
rect 267884 3380 267890 3392
rect 274818 3380 274824 3392
rect 267884 3352 274824 3380
rect 267884 3340 267890 3352
rect 274818 3340 274824 3352
rect 274876 3340 274882 3392
rect 300854 3340 300860 3392
rect 300912 3380 300918 3392
rect 310238 3380 310244 3392
rect 300912 3352 310244 3380
rect 300912 3340 300918 3352
rect 310238 3340 310244 3352
rect 310296 3340 310302 3392
rect 313366 3340 313372 3392
rect 313424 3380 313430 3392
rect 323302 3380 323308 3392
rect 313424 3352 323308 3380
rect 313424 3340 313430 3352
rect 323302 3340 323308 3352
rect 323360 3340 323366 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 352834 3380 352840 3392
rect 340932 3352 352840 3380
rect 340932 3340 340938 3352
rect 352834 3340 352840 3352
rect 352892 3340 352898 3392
rect 353294 3340 353300 3392
rect 353352 3380 353358 3392
rect 367002 3380 367008 3392
rect 353352 3352 367008 3380
rect 353352 3340 353358 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 378134 3340 378140 3392
rect 378192 3380 378198 3392
rect 393038 3380 393044 3392
rect 378192 3352 393044 3380
rect 378192 3340 378198 3352
rect 393038 3340 393044 3352
rect 393096 3340 393102 3392
rect 393314 3340 393320 3392
rect 393372 3380 393378 3392
rect 405016 3380 405044 3556
rect 410794 3544 410800 3556
rect 410852 3544 410858 3596
rect 411254 3544 411260 3596
rect 411312 3584 411318 3596
rect 429654 3584 429660 3596
rect 411312 3556 429660 3584
rect 411312 3544 411318 3556
rect 429654 3544 429660 3556
rect 429712 3544 429718 3596
rect 431926 3556 441614 3584
rect 407114 3476 407120 3528
rect 407172 3516 407178 3528
rect 424962 3516 424968 3528
rect 407172 3488 424968 3516
rect 407172 3476 407178 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 427814 3476 427820 3528
rect 427872 3516 427878 3528
rect 431926 3516 431954 3556
rect 427872 3488 431954 3516
rect 441586 3516 441614 3556
rect 442994 3544 443000 3596
rect 443052 3584 443058 3596
rect 463970 3584 463976 3596
rect 443052 3556 463976 3584
rect 443052 3544 443058 3556
rect 463970 3544 463976 3556
rect 464028 3544 464034 3596
rect 464338 3544 464344 3596
rect 464396 3584 464402 3596
rect 465166 3584 465172 3596
rect 464396 3556 465172 3584
rect 464396 3544 464402 3556
rect 465166 3544 465172 3556
rect 465224 3544 465230 3596
rect 470594 3544 470600 3596
rect 470652 3584 470658 3596
rect 493502 3584 493508 3596
rect 470652 3556 493508 3584
rect 470652 3544 470658 3556
rect 493502 3544 493508 3556
rect 493560 3544 493566 3596
rect 496814 3544 496820 3596
rect 496872 3584 496878 3596
rect 521838 3584 521844 3596
rect 496872 3556 521844 3584
rect 496872 3544 496878 3556
rect 521838 3544 521844 3556
rect 521896 3544 521902 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 539594 3584 539600 3596
rect 525116 3556 539600 3584
rect 525116 3544 525122 3556
rect 539594 3544 539600 3556
rect 539652 3544 539658 3596
rect 546494 3544 546500 3596
rect 546552 3584 546558 3596
rect 575106 3584 575112 3596
rect 546552 3556 575112 3584
rect 546552 3544 546558 3556
rect 575106 3544 575112 3556
rect 575164 3544 575170 3596
rect 447410 3516 447416 3528
rect 441586 3488 447416 3516
rect 427872 3476 427878 3488
rect 447410 3476 447416 3488
rect 447468 3476 447474 3528
rect 454678 3476 454684 3528
rect 454736 3516 454742 3528
rect 458082 3516 458088 3528
rect 454736 3488 458088 3516
rect 454736 3476 454742 3488
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 458192 3488 475332 3516
rect 417878 3448 417884 3460
rect 393372 3352 405044 3380
rect 408466 3420 417884 3448
rect 393372 3340 393378 3352
rect 20622 3272 20628 3324
rect 20680 3312 20686 3324
rect 25498 3312 25504 3324
rect 20680 3284 25504 3312
rect 20680 3272 20686 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 223666 3272 223672 3324
rect 223724 3312 223730 3324
rect 226334 3312 226340 3324
rect 223724 3284 226340 3312
rect 223724 3272 223730 3284
rect 226334 3272 226340 3284
rect 226392 3272 226398 3324
rect 238754 3272 238760 3324
rect 238812 3312 238818 3324
rect 242894 3312 242900 3324
rect 238812 3284 242900 3312
rect 238812 3272 238818 3284
rect 242894 3272 242900 3284
rect 242952 3272 242958 3324
rect 253934 3272 253940 3324
rect 253992 3312 253998 3324
rect 259454 3312 259460 3324
rect 253992 3284 259460 3312
rect 253992 3272 253998 3284
rect 259454 3272 259460 3284
rect 259512 3272 259518 3324
rect 296714 3272 296720 3324
rect 296772 3312 296778 3324
rect 305546 3312 305552 3324
rect 296772 3284 305552 3312
rect 296772 3272 296778 3284
rect 305546 3272 305552 3284
rect 305604 3272 305610 3324
rect 331214 3272 331220 3324
rect 331272 3312 331278 3324
rect 343358 3312 343364 3324
rect 331272 3284 343364 3312
rect 331272 3272 331278 3284
rect 343358 3272 343364 3284
rect 343416 3272 343422 3324
rect 345106 3272 345112 3324
rect 345164 3312 345170 3324
rect 358722 3312 358728 3324
rect 345164 3284 358728 3312
rect 345164 3272 345170 3284
rect 358722 3272 358728 3284
rect 358780 3272 358786 3324
rect 378226 3272 378232 3324
rect 378284 3312 378290 3324
rect 394234 3312 394240 3324
rect 378284 3284 394240 3312
rect 378284 3272 378290 3284
rect 394234 3272 394240 3284
rect 394292 3272 394298 3324
rect 402974 3272 402980 3324
rect 403032 3312 403038 3324
rect 407206 3312 407212 3324
rect 403032 3284 407212 3312
rect 403032 3272 403038 3284
rect 407206 3272 407212 3284
rect 407264 3272 407270 3324
rect 329926 3204 329932 3256
rect 329984 3244 329990 3256
rect 340966 3244 340972 3256
rect 329984 3216 340972 3244
rect 329984 3204 329990 3216
rect 340966 3204 340972 3216
rect 341024 3204 341030 3256
rect 341058 3204 341064 3256
rect 341116 3244 341122 3256
rect 354030 3244 354036 3256
rect 341116 3216 354036 3244
rect 341116 3204 341122 3216
rect 354030 3204 354036 3216
rect 354088 3204 354094 3256
rect 400306 3204 400312 3256
rect 400364 3244 400370 3256
rect 408466 3244 408494 3420
rect 417878 3408 417884 3420
rect 417936 3408 417942 3460
rect 420914 3408 420920 3460
rect 420972 3448 420978 3460
rect 420972 3420 438072 3448
rect 420972 3408 420978 3420
rect 411990 3340 411996 3392
rect 412048 3380 412054 3392
rect 422570 3380 422576 3392
rect 412048 3352 422576 3380
rect 412048 3340 412054 3352
rect 422570 3340 422576 3352
rect 422628 3340 422634 3392
rect 430942 3340 430948 3392
rect 431000 3380 431006 3392
rect 438044 3380 438072 3420
rect 438118 3408 438124 3460
rect 438176 3448 438182 3460
rect 439130 3448 439136 3460
rect 438176 3420 439136 3448
rect 438176 3408 438182 3420
rect 439130 3408 439136 3420
rect 439188 3408 439194 3460
rect 440326 3380 440332 3392
rect 431000 3352 431954 3380
rect 438044 3352 440332 3380
rect 431000 3340 431006 3352
rect 431926 3312 431954 3352
rect 440326 3340 440332 3352
rect 440384 3340 440390 3392
rect 449802 3380 449808 3392
rect 441586 3352 449808 3380
rect 441586 3312 441614 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 454034 3340 454040 3392
rect 454092 3380 454098 3392
rect 458192 3380 458220 3488
rect 458266 3408 458272 3460
rect 458324 3448 458330 3460
rect 475304 3448 475332 3488
rect 475378 3476 475384 3528
rect 475436 3516 475442 3528
rect 476942 3516 476948 3528
rect 475436 3488 476948 3516
rect 475436 3476 475442 3488
rect 476942 3476 476948 3488
rect 477000 3476 477006 3528
rect 478230 3476 478236 3528
rect 478288 3516 478294 3528
rect 485222 3516 485228 3528
rect 478288 3488 485228 3516
rect 478288 3476 478294 3488
rect 485222 3476 485228 3488
rect 485280 3476 485286 3528
rect 485774 3476 485780 3528
rect 485832 3516 485838 3528
rect 510062 3516 510068 3528
rect 485832 3488 510068 3516
rect 485832 3476 485838 3488
rect 510062 3476 510068 3488
rect 510120 3476 510126 3528
rect 512086 3476 512092 3528
rect 512144 3516 512150 3528
rect 538398 3516 538404 3528
rect 512144 3488 538404 3516
rect 512144 3476 512150 3488
rect 538398 3476 538404 3488
rect 538456 3476 538462 3528
rect 545114 3476 545120 3528
rect 545172 3516 545178 3528
rect 573910 3516 573916 3528
rect 545172 3488 573916 3516
rect 545172 3476 545178 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 475746 3448 475752 3460
rect 458324 3420 475240 3448
rect 475304 3420 475752 3448
rect 458324 3408 458330 3420
rect 472250 3380 472256 3392
rect 454092 3352 458220 3380
rect 460906 3352 472256 3380
rect 454092 3340 454098 3352
rect 431926 3284 441614 3312
rect 453298 3272 453304 3324
rect 453356 3312 453362 3324
rect 460906 3312 460934 3352
rect 472250 3340 472256 3352
rect 472308 3340 472314 3392
rect 475212 3380 475240 3420
rect 475746 3408 475752 3420
rect 475804 3408 475810 3460
rect 489914 3408 489920 3460
rect 489972 3448 489978 3460
rect 490742 3448 490748 3460
rect 489972 3420 490748 3448
rect 489972 3408 489978 3420
rect 490742 3408 490748 3420
rect 490800 3408 490806 3460
rect 514754 3448 514760 3460
rect 499546 3420 514760 3448
rect 479334 3380 479340 3392
rect 475212 3352 479340 3380
rect 479334 3340 479340 3352
rect 479392 3340 479398 3392
rect 490098 3340 490104 3392
rect 490156 3380 490162 3392
rect 499546 3380 499574 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 520274 3408 520280 3460
rect 520332 3448 520338 3460
rect 546678 3448 546684 3460
rect 520332 3420 546684 3448
rect 520332 3408 520338 3420
rect 546678 3408 546684 3420
rect 546736 3408 546742 3460
rect 553394 3408 553400 3460
rect 553452 3448 553458 3460
rect 583386 3448 583392 3460
rect 553452 3420 583392 3448
rect 553452 3408 553458 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 490156 3352 499574 3380
rect 490156 3340 490162 3352
rect 453356 3284 460934 3312
rect 453356 3272 453362 3284
rect 400364 3216 408494 3244
rect 400364 3204 400370 3216
rect 136450 3136 136456 3188
rect 136508 3176 136514 3188
rect 137278 3176 137284 3188
rect 136508 3148 137284 3176
rect 136508 3136 136514 3148
rect 137278 3136 137284 3148
rect 137336 3136 137342 3188
rect 201586 3136 201592 3188
rect 201644 3176 201650 3188
rect 203886 3176 203892 3188
rect 201644 3148 203892 3176
rect 201644 3136 201650 3148
rect 203886 3136 203892 3148
rect 203944 3136 203950 3188
rect 208670 3136 208676 3188
rect 208728 3176 208734 3188
rect 210970 3176 210976 3188
rect 208728 3148 210976 3176
rect 208728 3136 208734 3148
rect 210970 3136 210976 3148
rect 211028 3136 211034 3188
rect 215294 3136 215300 3188
rect 215352 3176 215358 3188
rect 218054 3176 218060 3188
rect 215352 3148 218060 3176
rect 215352 3136 215358 3148
rect 218054 3136 218060 3148
rect 218112 3136 218118 3188
rect 280154 3136 280160 3188
rect 280212 3176 280218 3188
rect 287790 3176 287796 3188
rect 280212 3148 287796 3176
rect 280212 3136 280218 3148
rect 287790 3136 287796 3148
rect 287848 3136 287854 3188
rect 324314 3136 324320 3188
rect 324372 3176 324378 3188
rect 335078 3176 335084 3188
rect 324372 3148 335084 3176
rect 324372 3136 324378 3148
rect 335078 3136 335084 3148
rect 335136 3136 335142 3188
rect 554038 3136 554044 3188
rect 554096 3176 554102 3188
rect 557350 3176 557356 3188
rect 554096 3148 557356 3176
rect 554096 3136 554102 3148
rect 557350 3136 557356 3148
rect 557408 3136 557414 3188
rect 255406 3068 255412 3120
rect 255464 3108 255470 3120
rect 260650 3108 260656 3120
rect 255464 3080 260656 3108
rect 255464 3068 255470 3080
rect 260650 3068 260656 3080
rect 260708 3068 260714 3120
rect 262214 3068 262220 3120
rect 262272 3108 262278 3120
rect 268838 3108 268844 3120
rect 262272 3080 268844 3108
rect 262272 3068 262278 3080
rect 268838 3068 268844 3080
rect 268896 3068 268902 3120
rect 278774 3068 278780 3120
rect 278832 3108 278838 3120
rect 286594 3108 286600 3120
rect 278832 3080 286600 3108
rect 278832 3068 278838 3080
rect 286594 3068 286600 3080
rect 286652 3068 286658 3120
rect 164878 3000 164884 3052
rect 164936 3040 164942 3052
rect 165706 3040 165712 3052
rect 164936 3012 165712 3040
rect 164936 3000 164942 3012
rect 165706 3000 165712 3012
rect 165764 3000 165770 3052
rect 167178 3000 167184 3052
rect 167236 3040 167242 3052
rect 168466 3040 168472 3052
rect 167236 3012 168472 3040
rect 167236 3000 167242 3012
rect 168466 3000 168472 3012
rect 168524 3000 168530 3052
rect 230474 3000 230480 3052
rect 230532 3040 230538 3052
rect 234614 3040 234620 3052
rect 230532 3012 234620 3040
rect 230532 3000 230538 3012
rect 234614 3000 234620 3012
rect 234672 3000 234678 3052
rect 289814 3000 289820 3052
rect 289872 3040 289878 3052
rect 298462 3040 298468 3052
rect 289872 3012 298468 3040
rect 289872 3000 289878 3012
rect 298462 3000 298468 3012
rect 298520 3000 298526 3052
rect 300118 3000 300124 3052
rect 300176 3040 300182 3052
rect 301958 3040 301964 3052
rect 300176 3012 301964 3040
rect 300176 3000 300182 3012
rect 301958 3000 301964 3012
rect 302016 3000 302022 3052
rect 476758 3000 476764 3052
rect 476816 3040 476822 3052
rect 481726 3040 481732 3052
rect 476816 3012 481732 3040
rect 476816 3000 476822 3012
rect 481726 3000 481732 3012
rect 481784 3000 481790 3052
rect 515398 3000 515404 3052
rect 515456 3040 515462 3052
rect 518342 3040 518348 3052
rect 515456 3012 518348 3040
rect 515456 3000 515462 3012
rect 518342 3000 518348 3012
rect 518400 3000 518406 3052
rect 73798 2932 73804 2984
rect 73856 2972 73862 2984
rect 75178 2972 75184 2984
rect 73856 2944 75184 2972
rect 73856 2932 73862 2944
rect 75178 2932 75184 2944
rect 75236 2932 75242 2984
rect 244366 2932 244372 2984
rect 244424 2972 244430 2984
rect 248782 2972 248788 2984
rect 244424 2944 248788 2972
rect 244424 2932 244430 2944
rect 248782 2932 248788 2944
rect 248840 2932 248846 2984
rect 281534 2932 281540 2984
rect 281592 2972 281598 2984
rect 288986 2972 288992 2984
rect 281592 2944 288992 2972
rect 281592 2932 281598 2944
rect 288986 2932 288992 2944
rect 289044 2932 289050 2984
rect 446398 2932 446404 2984
rect 446456 2972 446462 2984
rect 453298 2972 453304 2984
rect 446456 2944 453304 2972
rect 446456 2932 446462 2944
rect 453298 2932 453304 2944
rect 453356 2932 453362 2984
rect 287054 2864 287060 2916
rect 287112 2904 287118 2916
rect 296070 2904 296076 2916
rect 287112 2876 296076 2904
rect 287112 2864 287118 2876
rect 296070 2864 296076 2876
rect 296128 2864 296134 2916
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 218980 700884 219032 700936
rect 306380 700884 306432 700936
rect 264980 700816 265032 700868
rect 413652 700816 413704 700868
rect 154120 700748 154172 700800
rect 320180 700748 320232 700800
rect 137836 700680 137888 700732
rect 316040 700680 316092 700732
rect 249800 700612 249852 700664
rect 478512 700612 478564 700664
rect 89168 700544 89220 700596
rect 335360 700544 335412 700596
rect 72976 700476 73028 700528
rect 329840 700476 329892 700528
rect 236000 700408 236052 700460
rect 543464 700408 543516 700460
rect 24308 700340 24360 700392
rect 349160 700340 349212 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 218060 696940 218112 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 353944 683204 353996 683256
rect 222200 683136 222252 683188
rect 580172 683136 580224 683188
rect 282920 677220 282972 677272
rect 292856 677220 292908 677272
rect 278872 677152 278924 677204
rect 347780 677152 347832 677204
rect 269488 677084 269540 677136
rect 364340 677084 364392 677136
rect 201500 677016 201552 677068
rect 302240 677016 302292 677068
rect 255320 676948 255372 677000
rect 429200 676948 429252 677000
rect 241520 676880 241572 676932
rect 494060 676880 494112 676932
rect 227168 676812 227220 676864
rect 558920 676812 558972 676864
rect 266360 675724 266412 675776
rect 288440 675724 288492 675776
rect 274456 675656 274508 675708
rect 331220 675656 331272 675708
rect 260656 675588 260708 675640
rect 397460 675588 397512 675640
rect 246672 675520 246724 675572
rect 462320 675520 462372 675572
rect 232688 675452 232740 675504
rect 527180 675452 527232 675504
rect 194968 675384 195020 675436
rect 557172 675384 557224 675436
rect 180708 675316 180760 675368
rect 556988 675316 557040 675368
rect 166816 675248 166868 675300
rect 555976 675248 556028 675300
rect 157248 675180 157300 675232
rect 555884 675180 555936 675232
rect 148048 675112 148100 675164
rect 555792 675112 555844 675164
rect 133788 675044 133840 675096
rect 554596 675044 554648 675096
rect 119896 674976 119948 675028
rect 554412 674976 554464 675028
rect 91744 674908 91796 674960
rect 580172 674908 580224 674960
rect 4896 674840 4948 674892
rect 513748 674840 513800 674892
rect 284208 674364 284260 674416
rect 299480 674364 299532 674416
rect 234620 674296 234672 674348
rect 297732 674296 297784 674348
rect 169760 674228 169812 674280
rect 311900 674228 311952 674280
rect 104900 674160 104952 674212
rect 325884 674160 325936 674212
rect 40040 674092 40092 674144
rect 340052 674092 340104 674144
rect 204168 674024 204220 674076
rect 557356 674024 557408 674076
rect 13912 673956 13964 674008
rect 368572 673956 368624 674008
rect 8944 673888 8996 673940
rect 372804 673888 372856 673940
rect 11796 673820 11848 673872
rect 386972 673820 387024 673872
rect 6368 673752 6420 673804
rect 400956 673752 401008 673804
rect 6276 673684 6328 673736
rect 415492 673684 415544 673736
rect 6184 673616 6236 673668
rect 429200 673616 429252 673668
rect 5448 673548 5500 673600
rect 443276 673548 443328 673600
rect 3884 673480 3936 673532
rect 457444 673480 457496 673532
rect 198740 672936 198792 672988
rect 377588 672936 377640 672988
rect 175924 672868 175976 672920
rect 392032 672868 392084 672920
rect 395436 672868 395488 672920
rect 452660 672868 452712 672920
rect 105728 672800 105780 672852
rect 405740 672800 405792 672852
rect 115112 672732 115164 672784
rect 139492 672732 139544 672784
rect 152832 672732 152884 672784
rect 555700 672732 555752 672784
rect 10324 672664 10376 672716
rect 419724 672664 419776 672716
rect 419816 672664 419868 672716
rect 480812 672664 480864 672716
rect 138664 672596 138716 672648
rect 555608 672596 555660 672648
rect 13084 672528 13136 672580
rect 433892 672528 433944 672580
rect 54208 672460 54260 672512
rect 117964 672460 118016 672512
rect 124680 672460 124732 672512
rect 555516 672460 555568 672512
rect 4712 672392 4764 672444
rect 448060 672392 448112 672444
rect 448152 672392 448204 672444
rect 509240 672392 509292 672444
rect 5356 672324 5408 672376
rect 462320 672324 462372 672376
rect 96344 672256 96396 672308
rect 554136 672256 554188 672308
rect 5264 672188 5316 672240
rect 476212 672188 476264 672240
rect 5172 672120 5224 672172
rect 490196 672120 490248 672172
rect 5080 672052 5132 672104
rect 504364 672052 504416 672104
rect 3332 671508 3384 671560
rect 175924 671508 175976 671560
rect 199752 671508 199804 671560
rect 557264 671508 557316 671560
rect 3240 671440 3292 671492
rect 363420 671440 363472 671492
rect 3056 671372 3108 671424
rect 198740 671372 198792 671424
rect 213736 671372 213788 671424
rect 579620 671372 579672 671424
rect 13360 671304 13412 671356
rect 382280 671304 382332 671356
rect 397092 671304 397144 671356
rect 580540 671304 580592 671356
rect 185584 671236 185636 671288
rect 556068 671236 556120 671288
rect 176200 671168 176252 671220
rect 557080 671168 557132 671220
rect 171600 671100 171652 671152
rect 556896 671100 556948 671152
rect 13268 671032 13320 671084
rect 410340 671032 410392 671084
rect 13176 670964 13228 671016
rect 424508 670964 424560 671016
rect 129280 670896 129332 670948
rect 554504 670896 554556 670948
rect 3792 670828 3844 670880
rect 466828 670828 466880 670880
rect 72976 670760 73028 670812
rect 554044 670760 554096 670812
rect 3424 670692 3476 670744
rect 494980 670692 495032 670744
rect 3976 670216 4028 670268
rect 395436 670216 395488 670268
rect 209136 670148 209188 670200
rect 555332 670148 555384 670200
rect 3608 670080 3660 670132
rect 419816 670080 419868 670132
rect 190184 670012 190236 670064
rect 553952 670012 554004 670064
rect 4068 669944 4120 669996
rect 105728 669944 105780 669996
rect 117964 669944 118016 669996
rect 580356 669944 580408 669996
rect 143448 669876 143500 669928
rect 554688 669876 554740 669928
rect 110328 669808 110380 669860
rect 554228 669808 554280 669860
rect 105728 669740 105780 669792
rect 554320 669740 554372 669792
rect 86868 669672 86920 669724
rect 580908 669672 580960 669724
rect 58808 669604 58860 669656
rect 555424 669604 555476 669656
rect 82360 669536 82412 669588
rect 580724 669536 580776 669588
rect 77576 669468 77628 669520
rect 580816 669468 580868 669520
rect 63408 669400 63460 669452
rect 580632 669400 580684 669452
rect 49424 669332 49476 669384
rect 580448 669332 580500 669384
rect 3148 658180 3200 658232
rect 6460 658180 6512 658232
rect 557356 644376 557408 644428
rect 579988 644376 580040 644428
rect 3148 633360 3200 633412
rect 13820 633360 13872 633412
rect 555332 632000 555384 632052
rect 579988 632000 580040 632052
rect 557264 618196 557316 618248
rect 579988 618196 580040 618248
rect 3148 606772 3200 606824
rect 8944 606772 8996 606824
rect 553952 591948 554004 592000
rect 579804 591948 579856 592000
rect 3240 580932 3292 580984
rect 13360 580932 13412 580984
rect 557172 578144 557224 578196
rect 579804 578144 579856 578196
rect 556068 564340 556120 564392
rect 579988 564340 580040 564392
rect 3332 554684 3384 554736
rect 11796 554684 11848 554736
rect 557080 538160 557132 538212
rect 579988 538160 580040 538212
rect 556988 525716 557040 525768
rect 579988 525716 580040 525768
rect 556896 511912 556948 511964
rect 579988 511912 580040 511964
rect 3240 502120 3292 502172
rect 6368 502120 6420 502172
rect 3332 476008 3384 476060
rect 13268 476008 13320 476060
rect 555976 471928 556028 471980
rect 579804 471928 579856 471980
rect 3332 463632 3384 463684
rect 10324 463632 10376 463684
rect 555884 458124 555936 458176
rect 579988 458124 580040 458176
rect 3148 449556 3200 449608
rect 6276 449556 6328 449608
rect 555792 431876 555844 431928
rect 579988 431876 580040 431928
rect 3332 423580 3384 423632
rect 13176 423580 13228 423632
rect 555700 419432 555752 419484
rect 579988 419432 580040 419484
rect 3332 411204 3384 411256
rect 13084 411204 13136 411256
rect 554688 405628 554740 405680
rect 579988 405628 580040 405680
rect 3148 398692 3200 398744
rect 6184 398692 6236 398744
rect 554596 379448 554648 379500
rect 579804 379448 579856 379500
rect 555608 365644 555660 365696
rect 579988 365644 580040 365696
rect 2780 358436 2832 358488
rect 4712 358436 4764 358488
rect 554504 353200 554556 353252
rect 579988 353200 580040 353252
rect 2780 345856 2832 345908
rect 5448 345856 5500 345908
rect 554412 325592 554464 325644
rect 579988 325592 580040 325644
rect 555516 313216 555568 313268
rect 579988 313216 580040 313268
rect 2780 306212 2832 306264
rect 5356 306212 5408 306264
rect 554320 273164 554372 273216
rect 580080 273164 580132 273216
rect 554228 259360 554280 259412
rect 580080 259360 580132 259412
rect 2780 254328 2832 254380
rect 5264 254328 5316 254380
rect 556804 245556 556856 245608
rect 580080 245556 580132 245608
rect 554136 219376 554188 219428
rect 580172 219376 580224 219428
rect 2780 202376 2832 202428
rect 5172 202376 5224 202428
rect 554044 166948 554096 167000
rect 579620 166948 579672 167000
rect 2780 149880 2832 149932
rect 5080 149880 5132 149932
rect 3240 137912 3292 137964
rect 11704 137912 11756 137964
rect 555424 126896 555476 126948
rect 579620 126896 579672 126948
rect 2780 97860 2832 97912
rect 4988 97860 5040 97912
rect 2780 84872 2832 84924
rect 4896 84872 4948 84924
rect 2780 58624 2832 58676
rect 4804 58624 4856 58676
rect 22284 48220 22336 48272
rect 34980 48220 35032 48272
rect 35992 48220 36044 48272
rect 46940 48220 46992 48272
rect 55312 48220 55364 48272
rect 65524 48220 65576 48272
rect 68284 48220 68336 48272
rect 75460 48220 75512 48272
rect 100944 48220 100996 48272
rect 107292 48220 107344 48272
rect 434352 48220 434404 48272
rect 446404 48220 446456 48272
rect 463608 48220 463660 48272
rect 478052 48220 478104 48272
rect 11060 48152 11112 48204
rect 23940 48152 23992 48204
rect 24952 48152 25004 48204
rect 37280 48152 37332 48204
rect 41512 48152 41564 48204
rect 52460 48152 52512 48204
rect 52552 48152 52604 48204
rect 62212 48152 62264 48204
rect 96620 48152 96672 48204
rect 103980 48152 104032 48204
rect 416688 48152 416740 48204
rect 433340 48152 433392 48204
rect 438584 48152 438636 48204
rect 454684 48152 454736 48204
rect 460572 48152 460624 48204
rect 476764 48152 476816 48204
rect 478144 48152 478196 48204
rect 485044 48152 485096 48204
rect 514208 48152 514260 48204
rect 525064 48152 525116 48204
rect 16580 48084 16632 48136
rect 29460 48084 29512 48136
rect 44364 48084 44416 48136
rect 55772 48084 55824 48136
rect 60832 48084 60884 48136
rect 71044 48084 71096 48136
rect 199936 48084 199988 48136
rect 200120 48084 200172 48136
rect 409880 48084 409932 48136
rect 426440 48084 426492 48136
rect 433248 48084 433300 48136
rect 451280 48084 451332 48136
rect 469128 48084 469180 48136
rect 489920 48084 489972 48136
rect 494520 48084 494572 48136
rect 515404 48084 515456 48136
rect 530768 48084 530820 48136
rect 554044 48084 554096 48136
rect 15200 48016 15252 48068
rect 28356 48016 28408 48068
rect 38752 48016 38804 48068
rect 50252 48016 50304 48068
rect 56692 48016 56744 48068
rect 66628 48016 66680 48068
rect 69112 48016 69164 48068
rect 77668 48016 77720 48068
rect 80244 48016 80296 48068
rect 88524 48016 88576 48068
rect 91100 48016 91152 48068
rect 98460 48016 98512 48068
rect 103520 48016 103572 48068
rect 110420 48016 110472 48068
rect 111984 48016 112036 48068
rect 118148 48016 118200 48068
rect 414112 48016 414164 48068
rect 432144 48016 432196 48068
rect 446312 48016 446364 48068
rect 465264 48016 465316 48068
rect 474648 48016 474700 48068
rect 482284 48016 482336 48068
rect 11152 47948 11204 48000
rect 25044 47948 25096 48000
rect 31944 47948 31996 48000
rect 43628 47948 43680 48000
rect 51172 47948 51224 48000
rect 61108 47948 61160 48000
rect 63684 47948 63736 48000
rect 73252 47948 73304 48000
rect 78772 47948 78824 48000
rect 87420 47948 87472 48000
rect 89812 47948 89864 48000
rect 97356 47948 97408 48000
rect 104900 47948 104952 48000
rect 111800 47948 111852 48000
rect 113180 47948 113232 48000
rect 119252 47948 119304 48000
rect 420000 47948 420052 48000
rect 437480 47948 437532 48000
rect 439688 47948 439740 48000
rect 458180 47948 458232 48000
rect 462688 47948 462740 48000
rect 483020 48016 483072 48068
rect 488632 48016 488684 48068
rect 512000 48016 512052 48068
rect 515312 48016 515364 48068
rect 539784 48016 539836 48068
rect 483204 47948 483256 48000
rect 506664 47948 506716 48000
rect 508688 47948 508740 48000
rect 532700 47948 532752 48000
rect 537208 47948 537260 48000
rect 555424 48016 555476 48068
rect 550456 47948 550508 48000
rect 556896 47948 556948 48000
rect 12440 47880 12492 47932
rect 26332 47880 26384 47932
rect 33232 47880 33284 47932
rect 44732 47880 44784 47932
rect 45652 47880 45704 47932
rect 56876 47880 56928 47932
rect 59544 47880 59596 47932
rect 69020 47880 69072 47932
rect 71872 47880 71924 47932
rect 80980 47880 81032 47932
rect 92480 47880 92532 47932
rect 99564 47880 99616 47932
rect 109132 47880 109184 47932
rect 114836 47880 114888 47932
rect 127072 47880 127124 47932
rect 132592 47880 132644 47932
rect 144920 47880 144972 47932
rect 149060 47880 149112 47932
rect 151820 47880 151872 47932
rect 155316 47880 155368 47932
rect 161572 47880 161624 47932
rect 164240 47880 164292 47932
rect 230388 47880 230440 47932
rect 233240 47880 233292 47932
rect 372896 47880 372948 47932
rect 385684 47880 385736 47932
rect 393320 47880 393372 47932
rect 408500 47880 408552 47932
rect 423312 47880 423364 47932
rect 440424 47880 440476 47932
rect 445208 47880 445260 47932
rect 464344 47880 464396 47932
rect 466000 47880 466052 47932
rect 481272 47880 481324 47932
rect 482560 47880 482612 47932
rect 2780 47812 2832 47864
rect 17316 47812 17368 47864
rect 19616 47812 19668 47864
rect 31760 47812 31812 47864
rect 40132 47812 40184 47864
rect 51356 47812 51408 47864
rect 54024 47812 54076 47864
rect 64420 47812 64472 47864
rect 67824 47812 67876 47864
rect 76564 47812 76616 47864
rect 85764 47812 85816 47864
rect 94044 47812 94096 47864
rect 98092 47812 98144 47864
rect 105084 47812 105136 47864
rect 105544 47812 105596 47864
rect 108212 47812 108264 47864
rect 116032 47812 116084 47864
rect 121552 47812 121604 47864
rect 125600 47812 125652 47864
rect 130292 47812 130344 47864
rect 130476 47812 130528 47864
rect 131396 47812 131448 47864
rect 133880 47812 133932 47864
rect 138020 47812 138072 47864
rect 143816 47812 143868 47864
rect 146668 47812 146720 47864
rect 153384 47812 153436 47864
rect 156420 47812 156472 47864
rect 157432 47812 157484 47864
rect 160192 47812 160244 47864
rect 186320 47812 186372 47864
rect 187148 47812 187200 47864
rect 201592 47812 201644 47864
rect 202420 47812 202472 47864
rect 211896 47812 211948 47864
rect 212540 47812 212592 47864
rect 213000 47812 213052 47864
rect 213920 47812 213972 47864
rect 226064 47812 226116 47864
rect 227720 47812 227772 47864
rect 229376 47812 229428 47864
rect 231860 47812 231912 47864
rect 244280 47812 244332 47864
rect 245292 47812 245344 47864
rect 255320 47812 255372 47864
rect 256148 47812 256200 47864
rect 262128 47812 262180 47864
rect 264244 47812 264296 47864
rect 271880 47812 271932 47864
rect 277400 47812 277452 47864
rect 287060 47812 287112 47864
rect 287980 47812 288032 47864
rect 308036 47812 308088 47864
rect 309784 47812 309836 47864
rect 313280 47812 313332 47864
rect 314292 47812 314344 47864
rect 320088 47812 320140 47864
rect 323584 47812 323636 47864
rect 329840 47812 329892 47864
rect 330668 47812 330720 47864
rect 370688 47812 370740 47864
rect 383660 47812 383712 47864
rect 387248 47812 387300 47864
rect 401600 47812 401652 47864
rect 405648 47812 405700 47864
rect 411904 47812 411956 47864
rect 413560 47812 413612 47864
rect 430580 47812 430632 47864
rect 436560 47812 436612 47864
rect 455420 47812 455472 47864
rect 456892 47812 456944 47864
rect 457812 47812 457864 47864
rect 8300 47744 8352 47796
rect 22192 47744 22244 47796
rect 23480 47744 23532 47796
rect 36084 47744 36136 47796
rect 46940 47744 46992 47796
rect 57980 47744 58032 47796
rect 60740 47744 60792 47796
rect 69940 47744 69992 47796
rect 70400 47744 70452 47796
rect 80060 47744 80112 47796
rect 86960 47744 87012 47796
rect 95240 47744 95292 47796
rect 99380 47744 99432 47796
rect 106280 47744 106332 47796
rect 107660 47744 107712 47796
rect 113732 47744 113784 47796
rect 114560 47744 114612 47796
rect 120356 47744 120408 47796
rect 121460 47744 121512 47796
rect 126980 47744 127032 47796
rect 136640 47744 136692 47796
rect 141148 47744 141200 47796
rect 146300 47744 146352 47796
rect 149980 47744 150032 47796
rect 173900 47744 173952 47796
rect 175280 47744 175332 47796
rect 377312 47744 377364 47796
rect 390744 47744 390796 47796
rect 400128 47744 400180 47796
rect 415584 47744 415636 47796
rect 437388 47744 437440 47796
rect 451740 47744 451792 47796
rect 451832 47744 451884 47796
rect 453304 47744 453356 47796
rect 456248 47744 456300 47796
rect 475384 47812 475436 47864
rect 481456 47812 481508 47864
rect 486424 47812 486476 47864
rect 492312 47880 492364 47932
rect 514852 47880 514904 47932
rect 517428 47880 517480 47932
rect 542360 47880 542412 47932
rect 543648 47880 543700 47932
rect 548156 47880 548208 47932
rect 548248 47880 548300 47932
rect 505100 47812 505152 47864
rect 525892 47812 525944 47864
rect 526812 47812 526864 47864
rect 459468 47744 459520 47796
rect 480260 47744 480312 47796
rect 485688 47744 485740 47796
rect 507860 47744 507912 47796
rect 525248 47744 525300 47796
rect 549168 47812 549220 47864
rect 551284 47812 551336 47864
rect 550640 47744 550692 47796
rect 552664 47812 552716 47864
rect 560944 47812 560996 47864
rect 566464 47744 566516 47796
rect 6920 47676 6972 47728
rect 20720 47676 20772 47728
rect 27620 47676 27672 47728
rect 40316 47676 40368 47728
rect 48412 47676 48464 47728
rect 59452 47676 59504 47728
rect 62120 47676 62172 47728
rect 72148 47676 72200 47728
rect 75920 47676 75972 47728
rect 84292 47676 84344 47728
rect 88340 47676 88392 47728
rect 96712 47676 96764 47728
rect 102324 47676 102376 47728
rect 109316 47676 109368 47728
rect 110604 47676 110656 47728
rect 115940 47676 115992 47728
rect 124312 47676 124364 47728
rect 129188 47676 129240 47728
rect 132592 47676 132644 47728
rect 136732 47676 136784 47728
rect 151912 47676 151964 47728
rect 154580 47676 154632 47728
rect 362868 47676 362920 47728
rect 375380 47676 375432 47728
rect 380624 47676 380676 47728
rect 394700 47676 394752 47728
rect 397000 47676 397052 47728
rect 412640 47676 412692 47728
rect 426348 47676 426400 47728
rect 444380 47676 444432 47728
rect 449624 47676 449676 47728
rect 469220 47676 469272 47728
rect 472624 47676 472676 47728
rect 494060 47676 494112 47728
rect 495256 47676 495308 47728
rect 518900 47676 518952 47728
rect 536104 47676 536156 47728
rect 563060 47676 563112 47728
rect 5540 47608 5592 47660
rect 19524 47608 19576 47660
rect 29000 47608 29052 47660
rect 41420 47608 41472 47660
rect 42800 47608 42852 47660
rect 53932 47608 53984 47660
rect 57980 47608 58032 47660
rect 67732 47608 67784 47660
rect 69020 47608 69072 47660
rect 78864 47608 78916 47660
rect 81440 47608 81492 47660
rect 89720 47608 89772 47660
rect 95240 47608 95292 47660
rect 102876 47608 102928 47660
rect 106280 47608 106332 47660
rect 112628 47608 112680 47660
rect 131212 47608 131264 47660
rect 135628 47608 135680 47660
rect 137284 47608 137336 47660
rect 140044 47608 140096 47660
rect 147772 47608 147824 47660
rect 151084 47608 151136 47660
rect 158812 47608 158864 47660
rect 160836 47608 160888 47660
rect 162952 47608 163004 47660
rect 165620 47608 165672 47660
rect 168380 47608 168432 47660
rect 169760 47608 169812 47660
rect 234620 47608 234672 47660
rect 237380 47608 237432 47660
rect 239956 47608 240008 47660
rect 240784 47608 240836 47660
rect 243728 47608 243780 47660
rect 246304 47608 246356 47660
rect 350632 47608 350684 47660
rect 362224 47608 362276 47660
rect 367100 47608 367152 47660
rect 380900 47608 380952 47660
rect 383476 47608 383528 47660
rect 399024 47608 399076 47660
rect 403624 47608 403676 47660
rect 419540 47608 419592 47660
rect 420736 47608 420788 47660
rect 438124 47608 438176 47660
rect 442908 47608 442960 47660
rect 462320 47608 462372 47660
rect 468208 47608 468260 47660
rect 490012 47608 490064 47660
rect 498936 47608 498988 47660
rect 523224 47608 523276 47660
rect 528284 47608 528336 47660
rect 554780 47608 554832 47660
rect 4160 47540 4212 47592
rect 18420 47540 18472 47592
rect 20720 47540 20772 47592
rect 33876 47540 33928 47592
rect 35900 47540 35952 47592
rect 48320 47540 48372 47592
rect 52460 47540 52512 47592
rect 63500 47540 63552 47592
rect 64880 47540 64932 47592
rect 74540 47540 74592 47592
rect 75184 47540 75236 47592
rect 82084 47540 82136 47592
rect 82820 47540 82872 47592
rect 91192 47540 91244 47592
rect 93952 47540 94004 47592
rect 101772 47540 101824 47592
rect 110512 47540 110564 47592
rect 117320 47540 117372 47592
rect 122840 47540 122892 47592
rect 128452 47540 128504 47592
rect 143632 47540 143684 47592
rect 147864 47540 147916 47592
rect 154580 47540 154632 47592
rect 157524 47540 157576 47592
rect 265624 47540 265676 47592
rect 270500 47540 270552 47592
rect 293868 47540 293920 47592
rect 300124 47540 300176 47592
rect 347688 47540 347740 47592
rect 358084 47540 358136 47592
rect 373816 47540 373868 47592
rect 387800 47540 387852 47592
rect 390376 47540 390428 47592
rect 405740 47540 405792 47592
rect 406936 47540 406988 47592
rect 423864 47540 423916 47592
rect 429936 47540 429988 47592
rect 448612 47540 448664 47592
rect 451740 47540 451792 47592
rect 457076 47540 457128 47592
rect 9680 47472 9732 47524
rect 22836 47472 22888 47524
rect 26240 47472 26292 47524
rect 38108 47472 38160 47524
rect 49700 47472 49752 47524
rect 60188 47472 60240 47524
rect 84292 47472 84344 47524
rect 91836 47472 91888 47524
rect 142160 47472 142212 47524
rect 145564 47472 145616 47524
rect 156052 47472 156104 47524
rect 158720 47472 158772 47524
rect 427728 47472 427780 47524
rect 439504 47472 439556 47524
rect 452476 47472 452528 47524
rect 473544 47540 473596 47592
rect 475936 47540 475988 47592
rect 498200 47540 498252 47592
rect 502248 47540 502300 47592
rect 525800 47540 525852 47592
rect 535000 47540 535052 47592
rect 561680 47540 561732 47592
rect 481272 47472 481324 47524
rect 487160 47472 487212 47524
rect 521476 47472 521528 47524
rect 548064 47472 548116 47524
rect 548156 47472 548208 47524
rect 556804 47472 556856 47524
rect 17960 47404 18012 47456
rect 30564 47404 30616 47456
rect 34520 47404 34572 47456
rect 45836 47404 45888 47456
rect 74540 47404 74592 47456
rect 83188 47404 83240 47456
rect 207480 47404 207532 47456
rect 208400 47404 208452 47456
rect 13912 47336 13964 47388
rect 27252 47336 27304 47388
rect 37280 47336 37332 47388
rect 49148 47336 49200 47388
rect 135444 47336 135496 47388
rect 138940 47336 138992 47388
rect 165620 47336 165672 47388
rect 167460 47336 167512 47388
rect 519728 47336 519780 47388
rect 522304 47336 522356 47388
rect 551560 47336 551612 47388
rect 558184 47336 558236 47388
rect 27712 47268 27764 47320
rect 39212 47268 39264 47320
rect 44272 47268 44324 47320
rect 54668 47268 54720 47320
rect 85580 47268 85632 47320
rect 92940 47268 92992 47320
rect 93860 47268 93912 47320
rect 100760 47268 100812 47320
rect 237104 47268 237156 47320
rect 240140 47268 240192 47320
rect 522948 47268 523000 47320
rect 529204 47268 529256 47320
rect 25504 47200 25556 47252
rect 32772 47200 32824 47252
rect 124864 47200 124916 47252
rect 125876 47200 125928 47252
rect 172520 47200 172572 47252
rect 174084 47200 174136 47252
rect 117320 47064 117372 47116
rect 122932 47064 122984 47116
rect 118792 46996 118844 47048
rect 124772 46996 124824 47048
rect 130384 46996 130436 47048
rect 133420 46996 133472 47048
rect 139492 46996 139544 47048
rect 143540 46996 143592 47048
rect 150532 46996 150584 47048
rect 153292 46996 153344 47048
rect 160100 46996 160152 47048
rect 163044 46996 163096 47048
rect 77300 46928 77352 46980
rect 86316 46928 86368 46980
rect 118884 46928 118936 46980
rect 123668 46928 123720 46980
rect 140872 46928 140924 46980
rect 144460 46928 144512 46980
rect 149244 46928 149296 46980
rect 152188 46928 152240 46980
rect 160284 46928 160336 46980
rect 161940 46928 161992 46980
rect 169760 46928 169812 46980
rect 171876 46928 171928 46980
rect 179420 46928 179472 46980
rect 180800 46928 180852 46980
rect 219348 46928 219400 46980
rect 220084 46928 220136 46980
rect 362040 46928 362092 46980
rect 366364 46928 366416 46980
rect 487896 46928 487948 46980
rect 490564 46928 490616 46980
rect 223580 46452 223632 46504
rect 224500 46452 224552 46504
rect 160100 11704 160152 11756
rect 161296 11704 161348 11756
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 516140 5448 516192 5500
rect 541992 5448 542044 5500
rect 525984 5380 526036 5432
rect 552664 5380 552716 5432
rect 517520 5312 517572 5364
rect 544384 5312 544436 5364
rect 531320 5244 531372 5296
rect 558552 5244 558604 5296
rect 473360 5176 473412 5228
rect 495900 5176 495952 5228
rect 505192 5176 505244 5228
rect 530124 5176 530176 5228
rect 531504 5176 531556 5228
rect 559748 5176 559800 5228
rect 469312 5108 469364 5160
rect 492312 5108 492364 5160
rect 509240 5108 509292 5160
rect 534908 5108 534960 5160
rect 542452 5108 542504 5160
rect 570328 5108 570380 5160
rect 488540 5040 488592 5092
rect 513564 5040 513616 5092
rect 528560 5040 528612 5092
rect 556160 5040 556212 5092
rect 478880 4972 478932 5024
rect 501788 4972 501840 5024
rect 502340 4972 502392 5024
rect 527824 4972 527876 5024
rect 538220 4972 538272 5024
rect 566832 4972 566884 5024
rect 466460 4904 466512 4956
rect 488816 4904 488868 4956
rect 495440 4904 495492 4956
rect 520740 4904 520792 4956
rect 536840 4904 536892 4956
rect 565636 4904 565688 4956
rect 476120 4836 476172 4888
rect 499396 4836 499448 4888
rect 505284 4836 505336 4888
rect 531320 4836 531372 4888
rect 540980 4836 541032 4888
rect 569132 4836 569184 4888
rect 440332 4768 440384 4820
rect 460388 4768 460440 4820
rect 478972 4768 479024 4820
rect 502984 4768 503036 4820
rect 510712 4768 510764 4820
rect 537208 4768 537260 4820
rect 543740 4768 543792 4820
rect 572720 4768 572772 4820
rect 77392 4088 77444 4140
rect 85764 4088 85816 4140
rect 252560 4088 252612 4140
rect 258264 4088 258316 4140
rect 292580 4088 292632 4140
rect 300768 4088 300820 4140
rect 302240 4088 302292 4140
rect 311440 4088 311492 4140
rect 313280 4088 313332 4140
rect 324412 4088 324464 4140
rect 339500 4088 339552 4140
rect 351644 4088 351696 4140
rect 356060 4088 356112 4140
rect 369400 4088 369452 4140
rect 380992 4088 381044 4140
rect 396540 4088 396592 4140
rect 398840 4088 398892 4140
rect 399116 4088 399168 4140
rect 401692 4088 401744 4140
rect 418988 4088 419040 4140
rect 447140 4088 447192 4140
rect 467472 4088 467524 4140
rect 485044 4088 485096 4140
rect 500592 4088 500644 4140
rect 523132 4088 523184 4140
rect 524328 4088 524380 4140
rect 555424 4088 555476 4140
rect 564440 4088 564492 4140
rect 226432 4020 226484 4072
rect 229836 4020 229888 4072
rect 234712 4020 234764 4072
rect 239312 4020 239364 4072
rect 271972 4020 272024 4072
rect 279516 4020 279568 4072
rect 295340 4020 295392 4072
rect 304356 4020 304408 4072
rect 309784 4020 309836 4072
rect 317328 4020 317380 4072
rect 322940 4020 322992 4072
rect 333888 4020 333940 4072
rect 333980 4020 334032 4072
rect 345756 4020 345808 4072
rect 347780 4020 347832 4072
rect 361120 4020 361172 4072
rect 362960 4020 363012 4072
rect 377680 4020 377732 4072
rect 387892 4020 387944 4072
rect 263600 3952 263652 4004
rect 270040 3952 270092 4004
rect 298100 3952 298152 4004
rect 306748 3952 306800 4004
rect 310520 3952 310572 4004
rect 320916 3952 320968 4004
rect 323584 3952 323636 4004
rect 330392 3952 330444 4004
rect 338120 3952 338172 4004
rect 350448 3952 350500 4004
rect 356244 3952 356296 4004
rect 370596 3952 370648 4004
rect 371240 3952 371292 4004
rect 385960 3952 386012 4004
rect 391940 4020 391992 4072
rect 408408 4020 408460 4072
rect 408592 4020 408644 4072
rect 426164 4020 426216 4072
rect 441620 4020 441672 4072
rect 456064 4020 456116 4072
rect 490564 4020 490616 4072
rect 511264 4020 511316 4072
rect 529204 4020 529256 4072
rect 549076 4020 549128 4072
rect 556804 4020 556856 4072
rect 571524 4020 571576 4072
rect 264244 3884 264296 3936
rect 267740 3884 267792 3936
rect 277492 3884 277544 3936
rect 285404 3884 285456 3936
rect 285680 3884 285732 3936
rect 293684 3884 293736 3936
rect 303620 3884 303672 3936
rect 312636 3884 312688 3936
rect 318800 3884 318852 3936
rect 329196 3884 329248 3936
rect 332600 3884 332652 3936
rect 344560 3884 344612 3936
rect 345020 3884 345072 3936
rect 357532 3884 357584 3936
rect 360200 3884 360252 3936
rect 374092 3884 374144 3936
rect 383752 3884 383804 3936
rect 403624 3952 403676 4004
rect 409972 3952 410024 4004
rect 428464 3952 428516 4004
rect 430764 3952 430816 4004
rect 450912 3952 450964 4004
rect 456984 3952 457036 4004
rect 478144 3952 478196 4004
rect 492680 3952 492732 4004
rect 517152 3952 517204 4004
rect 522304 3952 522356 4004
rect 545488 3952 545540 4004
rect 560944 3952 560996 4004
rect 582196 3952 582248 4004
rect 102232 3816 102284 3868
rect 105544 3816 105596 3868
rect 227812 3816 227864 3868
rect 231032 3816 231084 3868
rect 247040 3816 247092 3868
rect 252376 3816 252428 3868
rect 281632 3816 281684 3868
rect 290188 3816 290240 3868
rect 306380 3816 306432 3868
rect 316224 3816 316276 3868
rect 317420 3816 317472 3868
rect 328000 3816 328052 3868
rect 329840 3816 329892 3868
rect 342168 3816 342220 3868
rect 354680 3816 354732 3868
rect 368204 3816 368256 3868
rect 368480 3816 368532 3868
rect 383568 3816 383620 3868
rect 399116 3884 399168 3936
rect 415492 3884 415544 3936
rect 423680 3884 423732 3936
rect 442632 3884 442684 3936
rect 447232 3884 447284 3936
rect 468668 3884 468720 3936
rect 486424 3884 486476 3936
rect 504180 3884 504232 3936
rect 506572 3884 506624 3936
rect 532516 3884 532568 3936
rect 556896 3884 556948 3936
rect 578608 3884 578660 3936
rect 400128 3816 400180 3868
rect 416780 3816 416832 3868
rect 435548 3816 435600 3868
rect 452660 3816 452712 3868
rect 474556 3816 474608 3868
rect 499580 3816 499632 3868
rect 524236 3816 524288 3868
rect 524328 3816 524380 3868
rect 550272 3816 550324 3868
rect 551284 3816 551336 3868
rect 577412 3816 577464 3868
rect 121092 3748 121144 3800
rect 124864 3748 124916 3800
rect 256700 3748 256752 3800
rect 262956 3748 263008 3800
rect 282920 3748 282972 3800
rect 291384 3748 291436 3800
rect 299480 3748 299532 3800
rect 309048 3748 309100 3800
rect 311900 3748 311952 3800
rect 322112 3748 322164 3800
rect 328460 3748 328512 3800
rect 339868 3748 339920 3800
rect 343640 3748 343692 3800
rect 356336 3748 356388 3800
rect 357440 3748 357492 3800
rect 2872 3544 2924 3596
rect 15292 3544 15344 3596
rect 237472 3680 237524 3732
rect 241704 3680 241756 3732
rect 249984 3680 250036 3732
rect 255872 3680 255924 3732
rect 266360 3680 266412 3732
rect 272432 3680 272484 3732
rect 273260 3680 273312 3732
rect 280712 3680 280764 3732
rect 305000 3680 305052 3732
rect 315028 3680 315080 3732
rect 316040 3680 316092 3732
rect 326804 3680 326856 3732
rect 327080 3680 327132 3732
rect 338672 3680 338724 3732
rect 349160 3680 349212 3732
rect 362316 3680 362368 3732
rect 364340 3748 364392 3800
rect 378876 3748 378928 3800
rect 397460 3748 397512 3800
rect 414296 3748 414348 3800
rect 418160 3748 418212 3800
rect 436744 3748 436796 3800
rect 439504 3748 439556 3800
rect 446220 3748 446272 3800
rect 449900 3748 449952 3800
rect 471060 3748 471112 3800
rect 482284 3748 482336 3800
rect 497096 3748 497148 3800
rect 499764 3748 499816 3800
rect 525432 3748 525484 3800
rect 525892 3748 525944 3800
rect 553768 3748 553820 3800
rect 558184 3748 558236 3800
rect 581000 3748 581052 3800
rect 209780 3612 209832 3664
rect 212172 3612 212224 3664
rect 212632 3612 212684 3664
rect 215668 3612 215720 3664
rect 276020 3612 276072 3664
rect 283104 3612 283156 3664
rect 284300 3612 284352 3664
rect 292580 3612 292632 3664
rect 293960 3612 294012 3664
rect 303160 3612 303212 3664
rect 307760 3612 307812 3664
rect 318524 3612 318576 3664
rect 320180 3612 320232 3664
rect 331588 3612 331640 3664
rect 335360 3612 335412 3664
rect 346952 3612 347004 3664
rect 351920 3612 351972 3664
rect 365812 3612 365864 3664
rect 367192 3680 367244 3732
rect 382372 3680 382424 3732
rect 385040 3680 385092 3732
rect 401324 3680 401376 3732
rect 371700 3612 371752 3664
rect 375472 3612 375524 3664
rect 390560 3612 390612 3664
rect 390652 3612 390704 3664
rect 402980 3612 403032 3664
rect 16672 3544 16724 3596
rect 130568 3544 130620 3596
rect 133972 3544 134024 3596
rect 138848 3544 138900 3596
rect 142252 3544 142304 3596
rect 143632 3544 143684 3596
rect 144736 3544 144788 3596
rect 191932 3544 191984 3596
rect 193220 3544 193272 3596
rect 197452 3544 197504 3596
rect 199108 3544 199160 3596
rect 200212 3544 200264 3596
rect 201500 3544 201552 3596
rect 204352 3544 204404 3596
rect 206192 3544 206244 3596
rect 207020 3544 207072 3596
rect 1676 3476 1728 3528
rect 214012 3544 214064 3596
rect 216864 3544 216916 3596
rect 218060 3544 218112 3596
rect 220452 3544 220504 3596
rect 223580 3544 223632 3596
rect 227536 3544 227588 3596
rect 233332 3544 233384 3596
rect 237012 3544 237064 3596
rect 244280 3544 244332 3596
rect 249984 3544 250036 3596
rect 251180 3544 251232 3596
rect 257068 3544 257120 3596
rect 259460 3544 259512 3596
rect 265348 3544 265400 3596
rect 266452 3544 266504 3596
rect 273628 3544 273680 3596
rect 274640 3544 274692 3596
rect 281908 3544 281960 3596
rect 287152 3544 287204 3596
rect 294880 3544 294932 3596
rect 303712 3544 303764 3596
rect 313832 3544 313884 3596
rect 314660 3544 314712 3596
rect 325608 3544 325660 3596
rect 325700 3544 325752 3596
rect 337476 3544 337528 3596
rect 342260 3544 342312 3596
rect 355232 3544 355284 3596
rect 358820 3544 358872 3596
rect 372896 3544 372948 3596
rect 374000 3544 374052 3596
rect 389456 3544 389508 3596
rect 394792 3544 394844 3596
rect 411904 3680 411956 3732
rect 404360 3612 404412 3664
rect 421380 3680 421432 3732
rect 425060 3680 425112 3732
rect 443828 3680 443880 3732
rect 456064 3680 456116 3732
rect 461584 3680 461636 3732
rect 463700 3680 463752 3732
rect 486424 3680 486476 3732
rect 503720 3680 503772 3732
rect 529020 3680 529072 3732
rect 532792 3680 532844 3732
rect 560852 3680 560904 3732
rect 566464 3680 566516 3732
rect 576308 3680 576360 3732
rect 414020 3612 414072 3664
rect 433248 3612 433300 3664
rect 434720 3612 434772 3664
rect 454500 3612 454552 3664
rect 456800 3612 456852 3664
rect 458272 3612 458324 3664
rect 460940 3612 460992 3664
rect 482836 3612 482888 3664
rect 483112 3612 483164 3664
rect 507676 3612 507728 3664
rect 510620 3612 510672 3664
rect 536104 3612 536156 3664
rect 539692 3612 539744 3664
rect 568028 3612 568080 3664
rect 27620 3476 27672 3528
rect 28540 3476 28592 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 66720 3476 66772 3528
rect 68284 3476 68336 3528
rect 69020 3476 69072 3528
rect 69940 3476 69992 3528
rect 110512 3476 110564 3528
rect 111616 3476 111668 3528
rect 118792 3476 118844 3528
rect 119896 3476 119948 3528
rect 126980 3476 127032 3528
rect 128176 3476 128228 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 169760 3476 169812 3528
rect 170404 3476 170456 3528
rect 172520 3476 172572 3528
rect 172796 3476 172848 3528
rect 179052 3476 179104 3528
rect 179512 3476 179564 3528
rect 186320 3476 186372 3528
rect 186964 3476 187016 3528
rect 205640 3476 205692 3528
rect 207388 3476 207440 3528
rect 209780 3476 209832 3528
rect 216680 3476 216732 3528
rect 219256 3476 219308 3528
rect 220084 3476 220136 3528
rect 221556 3476 221608 3528
rect 222200 3476 222252 3528
rect 225144 3476 225196 3528
rect 231952 3476 232004 3528
rect 235816 3476 235868 3528
rect 240784 3476 240836 3528
rect 244096 3476 244148 3528
rect 246304 3476 246356 3528
rect 247592 3476 247644 3528
rect 249800 3476 249852 3528
rect 254676 3476 254728 3528
rect 255320 3476 255372 3528
rect 261760 3476 261812 3528
rect 270592 3476 270644 3528
rect 277124 3476 277176 3528
rect 291200 3476 291252 3528
rect 299664 3476 299716 3528
rect 309140 3476 309192 3528
rect 319720 3476 319772 3528
rect 321560 3476 321612 3528
rect 332692 3476 332744 3528
rect 335452 3476 335504 3528
rect 348056 3476 348108 3528
rect 350540 3476 350592 3528
rect 572 3408 624 3460
rect 13820 3408 13872 3460
rect 31300 3408 31352 3460
rect 42892 3408 42944 3460
rect 220820 3408 220872 3460
rect 223948 3408 224000 3460
rect 240232 3408 240284 3460
rect 245200 3408 245252 3460
rect 245660 3408 245712 3460
rect 251180 3408 251232 3460
rect 260840 3408 260892 3460
rect 266544 3408 266596 3460
rect 269120 3408 269172 3460
rect 276020 3408 276072 3460
rect 276112 3408 276164 3460
rect 284300 3408 284352 3460
rect 288440 3408 288492 3460
rect 297272 3408 297324 3460
rect 298192 3408 298244 3460
rect 307944 3408 307996 3460
rect 324504 3408 324556 3460
rect 336280 3408 336332 3460
rect 336740 3408 336792 3460
rect 349252 3408 349304 3460
rect 358084 3476 358136 3528
rect 359924 3476 359976 3528
rect 362224 3476 362276 3528
rect 363512 3476 363564 3528
rect 365720 3476 365772 3528
rect 379980 3476 380032 3528
rect 385684 3476 385736 3528
rect 387156 3476 387208 3528
rect 388076 3476 388128 3528
rect 404820 3476 404872 3528
rect 364616 3408 364668 3460
rect 366364 3408 366416 3460
rect 375288 3408 375340 3460
rect 382280 3408 382332 3460
rect 397736 3408 397788 3460
rect 126980 3340 127032 3392
rect 130476 3340 130528 3392
rect 219440 3340 219492 3392
rect 222752 3340 222804 3392
rect 241520 3340 241572 3392
rect 246396 3340 246448 3392
rect 248420 3340 248472 3392
rect 253480 3340 253532 3392
rect 258080 3340 258132 3392
rect 264152 3340 264204 3392
rect 267832 3340 267884 3392
rect 274824 3340 274876 3392
rect 300860 3340 300912 3392
rect 310244 3340 310296 3392
rect 313372 3340 313424 3392
rect 323308 3340 323360 3392
rect 340880 3340 340932 3392
rect 352840 3340 352892 3392
rect 353300 3340 353352 3392
rect 367008 3340 367060 3392
rect 378140 3340 378192 3392
rect 393044 3340 393096 3392
rect 393320 3340 393372 3392
rect 410800 3544 410852 3596
rect 411260 3544 411312 3596
rect 429660 3544 429712 3596
rect 407120 3476 407172 3528
rect 424968 3476 425020 3528
rect 427820 3476 427872 3528
rect 443000 3544 443052 3596
rect 463976 3544 464028 3596
rect 464344 3544 464396 3596
rect 465172 3544 465224 3596
rect 470600 3544 470652 3596
rect 493508 3544 493560 3596
rect 496820 3544 496872 3596
rect 521844 3544 521896 3596
rect 525064 3544 525116 3596
rect 539600 3544 539652 3596
rect 546500 3544 546552 3596
rect 575112 3544 575164 3596
rect 447416 3476 447468 3528
rect 454684 3476 454736 3528
rect 458088 3476 458140 3528
rect 20628 3272 20680 3324
rect 25504 3272 25556 3324
rect 223672 3272 223724 3324
rect 226340 3272 226392 3324
rect 238760 3272 238812 3324
rect 242900 3272 242952 3324
rect 253940 3272 253992 3324
rect 259460 3272 259512 3324
rect 296720 3272 296772 3324
rect 305552 3272 305604 3324
rect 331220 3272 331272 3324
rect 343364 3272 343416 3324
rect 345112 3272 345164 3324
rect 358728 3272 358780 3324
rect 378232 3272 378284 3324
rect 394240 3272 394292 3324
rect 402980 3272 403032 3324
rect 407212 3272 407264 3324
rect 329932 3204 329984 3256
rect 340972 3204 341024 3256
rect 341064 3204 341116 3256
rect 354036 3204 354088 3256
rect 400312 3204 400364 3256
rect 417884 3408 417936 3460
rect 420920 3408 420972 3460
rect 411996 3340 412048 3392
rect 422576 3340 422628 3392
rect 430948 3340 431000 3392
rect 438124 3408 438176 3460
rect 439136 3408 439188 3460
rect 440332 3340 440384 3392
rect 449808 3340 449860 3392
rect 454040 3340 454092 3392
rect 458272 3408 458324 3460
rect 475384 3476 475436 3528
rect 476948 3476 477000 3528
rect 478236 3476 478288 3528
rect 485228 3476 485280 3528
rect 485780 3476 485832 3528
rect 510068 3476 510120 3528
rect 512092 3476 512144 3528
rect 538404 3476 538456 3528
rect 545120 3476 545172 3528
rect 573916 3476 573968 3528
rect 453304 3272 453356 3324
rect 472256 3340 472308 3392
rect 475752 3408 475804 3460
rect 489920 3408 489972 3460
rect 490748 3408 490800 3460
rect 479340 3340 479392 3392
rect 490104 3340 490156 3392
rect 514760 3408 514812 3460
rect 520280 3408 520332 3460
rect 546684 3408 546736 3460
rect 553400 3408 553452 3460
rect 583392 3408 583444 3460
rect 136456 3136 136508 3188
rect 137284 3136 137336 3188
rect 201592 3136 201644 3188
rect 203892 3136 203944 3188
rect 208676 3136 208728 3188
rect 210976 3136 211028 3188
rect 215300 3136 215352 3188
rect 218060 3136 218112 3188
rect 280160 3136 280212 3188
rect 287796 3136 287848 3188
rect 324320 3136 324372 3188
rect 335084 3136 335136 3188
rect 554044 3136 554096 3188
rect 557356 3136 557408 3188
rect 255412 3068 255464 3120
rect 260656 3068 260708 3120
rect 262220 3068 262272 3120
rect 268844 3068 268896 3120
rect 278780 3068 278832 3120
rect 286600 3068 286652 3120
rect 164884 3000 164936 3052
rect 165712 3000 165764 3052
rect 167184 3000 167236 3052
rect 168472 3000 168524 3052
rect 230480 3000 230532 3052
rect 234620 3000 234672 3052
rect 289820 3000 289872 3052
rect 298468 3000 298520 3052
rect 300124 3000 300176 3052
rect 301964 3000 302016 3052
rect 476764 3000 476816 3052
rect 481732 3000 481784 3052
rect 515404 3000 515456 3052
rect 518348 3000 518400 3052
rect 73804 2932 73856 2984
rect 75184 2932 75236 2984
rect 244372 2932 244424 2984
rect 248788 2932 248840 2984
rect 281540 2932 281592 2984
rect 288992 2932 289044 2984
rect 446404 2932 446456 2984
rect 453304 2932 453356 2984
rect 287060 2864 287112 2916
rect 296076 2864 296128 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 4896 674892 4948 674898
rect 4896 674834 4948 674840
rect 3698 673840 3754 673849
rect 3698 673775 3754 673784
rect 3606 673704 3662 673713
rect 3606 673639 3662 673648
rect 3620 673454 3648 673639
rect 3528 673426 3648 673454
rect 3332 671560 3384 671566
rect 3332 671502 3384 671508
rect 3240 671492 3292 671498
rect 3240 671434 3292 671440
rect 3056 671424 3108 671430
rect 3056 671366 3108 671372
rect 3068 667298 3096 671366
rect 3252 671265 3280 671434
rect 3238 671256 3294 671265
rect 3238 671191 3294 671200
rect 3068 667270 3280 667298
rect 3148 658232 3200 658238
rect 3146 658200 3148 658209
rect 3200 658200 3202 658209
rect 3146 658135 3202 658144
rect 3148 633412 3200 633418
rect 3148 633354 3200 633360
rect 3160 632097 3188 633354
rect 3146 632088 3202 632097
rect 3146 632023 3202 632032
rect 3252 619177 3280 667270
rect 3238 619168 3294 619177
rect 3238 619103 3294 619112
rect 3148 606824 3200 606830
rect 3148 606766 3200 606772
rect 3160 606121 3188 606766
rect 3146 606112 3202 606121
rect 3146 606047 3202 606056
rect 3240 580984 3292 580990
rect 3240 580926 3292 580932
rect 3252 580009 3280 580926
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 671502
rect 3424 670744 3476 670750
rect 3424 670686 3476 670692
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3332 554736 3384 554742
rect 3332 554678 3384 554684
rect 3344 553897 3372 554678
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3240 502172 3292 502178
rect 3240 502114 3292 502120
rect 3252 501809 3280 502114
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3332 476060 3384 476066
rect 3332 476002 3384 476008
rect 3344 475697 3372 476002
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3332 463684 3384 463690
rect 3332 463626 3384 463632
rect 3344 462641 3372 463626
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3148 449608 3200 449614
rect 3146 449576 3148 449585
rect 3200 449576 3202 449585
rect 3146 449511 3202 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3148 398744 3200 398750
rect 3148 398686 3200 398692
rect 3160 397497 3188 398686
rect 3146 397488 3202 397497
rect 3146 397423 3202 397432
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 2780 345908 2832 345914
rect 2780 345850 2832 345856
rect 2792 345409 2820 345850
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2780 306264 2832 306270
rect 2778 306232 2780 306241
rect 2832 306232 2834 306241
rect 2778 306167 2834 306176
rect 2780 254380 2832 254386
rect 2780 254322 2832 254328
rect 2792 254153 2820 254322
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 2780 202428 2832 202434
rect 2780 202370 2832 202376
rect 2792 201929 2820 202370
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 3436 162897 3464 670686
rect 3528 188873 3556 673426
rect 3608 670132 3660 670138
rect 3608 670074 3660 670080
rect 3620 214985 3648 670074
rect 3712 241097 3740 673775
rect 3884 673532 3936 673538
rect 3884 673474 3936 673480
rect 3792 670880 3844 670886
rect 3792 670822 3844 670828
rect 3804 267209 3832 670822
rect 3896 293185 3924 673474
rect 4802 672616 4858 672625
rect 4802 672551 4858 672560
rect 4712 672444 4764 672450
rect 4712 672386 4764 672392
rect 3976 670268 4028 670274
rect 3976 670210 4028 670216
rect 3988 319297 4016 670210
rect 4068 669996 4120 670002
rect 4068 669938 4120 669944
rect 4080 514865 4108 669938
rect 4066 514856 4122 514865
rect 4066 514791 4122 514800
rect 4724 358494 4752 672386
rect 4712 358488 4764 358494
rect 4712 358430 4764 358436
rect 3974 319288 4030 319297
rect 3974 319223 4030 319232
rect 3882 293176 3938 293185
rect 3882 293111 3938 293120
rect 3790 267200 3846 267209
rect 3790 267135 3846 267144
rect 3698 241088 3754 241097
rect 3698 241023 3754 241032
rect 3606 214976 3662 214985
rect 3606 214911 3662 214920
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 2780 149932 2832 149938
rect 2780 149874 2832 149880
rect 2792 149841 2820 149874
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 2780 97912 2832 97918
rect 2780 97854 2832 97860
rect 2792 97617 2820 97854
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 2780 84924 2832 84930
rect 2780 84866 2832 84872
rect 2792 84697 2820 84866
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 4816 58682 4844 672551
rect 4908 84930 4936 674834
rect 40052 674150 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700534 73016 703520
rect 89180 700602 89208 703520
rect 89168 700596 89220 700602
rect 89168 700538 89220 700544
rect 72976 700528 73028 700534
rect 72976 700470 73028 700476
rect 91744 674960 91796 674966
rect 91744 674902 91796 674908
rect 40040 674144 40092 674150
rect 40040 674086 40092 674092
rect 13912 674008 13964 674014
rect 13912 673950 13964 673956
rect 8944 673940 8996 673946
rect 8944 673882 8996 673888
rect 6368 673804 6420 673810
rect 6368 673746 6420 673752
rect 6276 673736 6328 673742
rect 6276 673678 6328 673684
rect 6184 673668 6236 673674
rect 6184 673610 6236 673616
rect 5448 673600 5500 673606
rect 5448 673542 5500 673548
rect 5356 672376 5408 672382
rect 4986 672344 5042 672353
rect 5356 672318 5408 672324
rect 4986 672279 5042 672288
rect 5000 97918 5028 672279
rect 5264 672240 5316 672246
rect 5264 672182 5316 672188
rect 5172 672172 5224 672178
rect 5172 672114 5224 672120
rect 5080 672104 5132 672110
rect 5080 672046 5132 672052
rect 5092 149938 5120 672046
rect 5184 202434 5212 672114
rect 5276 254386 5304 672182
rect 5368 306270 5396 672318
rect 5460 345914 5488 673542
rect 6196 398750 6224 673610
rect 6288 449614 6316 673678
rect 6380 502178 6408 673746
rect 6458 668128 6514 668137
rect 6458 668063 6514 668072
rect 6472 658238 6500 668063
rect 6460 658232 6512 658238
rect 6460 658174 6512 658180
rect 8956 606830 8984 673882
rect 11796 673872 11848 673878
rect 11796 673814 11848 673820
rect 11702 673568 11758 673577
rect 11702 673503 11758 673512
rect 10324 672716 10376 672722
rect 10324 672658 10376 672664
rect 8944 606824 8996 606830
rect 8944 606766 8996 606772
rect 6368 502172 6420 502178
rect 6368 502114 6420 502120
rect 10336 463690 10364 672658
rect 10324 463684 10376 463690
rect 10324 463626 10376 463632
rect 6276 449608 6328 449614
rect 6276 449550 6328 449556
rect 6184 398744 6236 398750
rect 6184 398686 6236 398692
rect 5448 345908 5500 345914
rect 5448 345850 5500 345856
rect 5356 306264 5408 306270
rect 5356 306206 5408 306212
rect 5264 254380 5316 254386
rect 5264 254322 5316 254328
rect 5172 202428 5224 202434
rect 5172 202370 5224 202376
rect 5080 149932 5132 149938
rect 5080 149874 5132 149880
rect 11716 137970 11744 673503
rect 11808 554742 11836 673814
rect 13084 672580 13136 672586
rect 13084 672522 13136 672528
rect 11796 554736 11848 554742
rect 11796 554678 11848 554684
rect 13096 411262 13124 672522
rect 13360 671356 13412 671362
rect 13360 671298 13412 671304
rect 13268 671084 13320 671090
rect 13268 671026 13320 671032
rect 13176 671016 13228 671022
rect 13176 670958 13228 670964
rect 13188 423638 13216 670958
rect 13280 476066 13308 671026
rect 13372 580990 13400 671298
rect 13924 634814 13952 673950
rect 54208 672512 54260 672518
rect 54208 672454 54260 672460
rect 68190 672480 68246 672489
rect 44822 670848 44878 670857
rect 44822 670783 44878 670792
rect 44836 669882 44864 670783
rect 54220 669882 54248 672454
rect 68190 672415 68246 672424
rect 68204 669882 68232 672415
rect 72976 670812 73028 670818
rect 72976 670754 73028 670760
rect 72988 669882 73016 670754
rect 91756 669882 91784 674902
rect 104912 674218 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 700738 137876 703520
rect 154132 700806 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700800 154172 700806
rect 154120 700742 154172 700748
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 166816 675300 166868 675306
rect 166816 675242 166868 675248
rect 157248 675232 157300 675238
rect 157248 675174 157300 675180
rect 148048 675164 148100 675170
rect 148048 675106 148100 675112
rect 133788 675096 133840 675102
rect 133788 675038 133840 675044
rect 119896 675028 119948 675034
rect 119896 674970 119948 674976
rect 104900 674212 104952 674218
rect 104900 674154 104952 674160
rect 101126 673976 101182 673985
rect 101126 673911 101182 673920
rect 96344 672308 96396 672314
rect 96344 672250 96396 672256
rect 96356 669882 96384 672250
rect 101140 669882 101168 673911
rect 105728 672852 105780 672858
rect 105728 672794 105780 672800
rect 105740 670002 105768 672794
rect 115112 672784 115164 672790
rect 115112 672726 115164 672732
rect 105728 669996 105780 670002
rect 105728 669938 105780 669944
rect 115124 669882 115152 672726
rect 117964 672512 118016 672518
rect 117964 672454 118016 672460
rect 117976 670002 118004 672454
rect 117964 669996 118016 670002
rect 117964 669938 118016 669944
rect 119908 669882 119936 674970
rect 124680 672512 124732 672518
rect 124680 672454 124732 672460
rect 124692 669882 124720 672454
rect 129280 670948 129332 670954
rect 129280 670890 129332 670896
rect 129292 669882 129320 670890
rect 133800 669882 133828 675038
rect 139492 672784 139544 672790
rect 139492 672726 139544 672732
rect 138664 672648 138716 672654
rect 138664 672590 138716 672596
rect 138676 669882 138704 672590
rect 44482 669854 44864 669882
rect 53866 669854 54248 669882
rect 67942 669854 68232 669882
rect 72634 669854 73016 669882
rect 91402 669854 91784 669882
rect 96094 669854 96384 669882
rect 100786 669854 101168 669882
rect 110170 669866 110368 669882
rect 110170 669860 110380 669866
rect 110170 669854 110328 669860
rect 114862 669854 115152 669882
rect 119554 669854 119936 669882
rect 124338 669854 124720 669882
rect 129030 669854 129320 669882
rect 133722 669854 133828 669882
rect 138414 669854 138704 669882
rect 110328 669802 110380 669808
rect 105728 669792 105780 669798
rect 86710 669730 86908 669746
rect 105478 669740 105728 669746
rect 105478 669734 105780 669740
rect 86710 669724 86920 669730
rect 86710 669718 86868 669724
rect 105478 669718 105768 669734
rect 86868 669666 86920 669672
rect 58808 669656 58860 669662
rect 58558 669604 58808 669610
rect 139504 669633 139532 672726
rect 143448 669928 143500 669934
rect 143106 669876 143448 669882
rect 148060 669882 148088 675106
rect 152832 672784 152884 672790
rect 152832 672726 152884 672732
rect 152844 669882 152872 672726
rect 157260 669882 157288 675174
rect 166828 669882 166856 675242
rect 169772 674286 169800 702406
rect 201512 677074 201540 702986
rect 218992 700942 219020 703520
rect 218980 700936 219032 700942
rect 218980 700878 219032 700884
rect 218060 696992 218112 696998
rect 218060 696934 218112 696940
rect 201500 677068 201552 677074
rect 201500 677010 201552 677016
rect 194968 675436 195020 675442
rect 194968 675378 195020 675384
rect 180708 675368 180760 675374
rect 180708 675310 180760 675316
rect 169760 674280 169812 674286
rect 169760 674222 169812 674228
rect 175924 672920 175976 672926
rect 175924 672862 175976 672868
rect 175936 671566 175964 672862
rect 175924 671560 175976 671566
rect 175924 671502 175976 671508
rect 176200 671220 176252 671226
rect 176200 671162 176252 671168
rect 171600 671152 171652 671158
rect 171600 671094 171652 671100
rect 171612 669882 171640 671094
rect 176212 669882 176240 671162
rect 180720 669882 180748 675310
rect 185584 671288 185636 671294
rect 185584 671230 185636 671236
rect 185596 669882 185624 671230
rect 190184 670064 190236 670070
rect 190184 670006 190236 670012
rect 190196 669882 190224 670006
rect 194980 669882 195008 675378
rect 204168 674076 204220 674082
rect 204168 674018 204220 674024
rect 198740 672988 198792 672994
rect 198740 672930 198792 672936
rect 198752 671430 198780 672930
rect 199752 671560 199804 671566
rect 199752 671502 199804 671508
rect 198740 671424 198792 671430
rect 198740 671366 198792 671372
rect 199764 669882 199792 671502
rect 204180 669882 204208 674018
rect 213736 671424 213788 671430
rect 213736 671366 213788 671372
rect 209136 670200 209188 670206
rect 209136 670142 209188 670148
rect 209148 669882 209176 670142
rect 213748 669882 213776 671366
rect 143106 669870 143500 669876
rect 143106 669854 143488 669870
rect 147798 669854 148088 669882
rect 152490 669854 152872 669882
rect 157182 669854 157288 669882
rect 166566 669854 166856 669882
rect 171258 669854 171640 669882
rect 175950 669854 176240 669882
rect 180642 669854 180748 669882
rect 185334 669854 185624 669882
rect 190026 669854 190224 669882
rect 194718 669854 195008 669882
rect 199410 669854 199792 669882
rect 204102 669854 204208 669882
rect 208794 669854 209176 669882
rect 213486 669854 213776 669882
rect 218072 669882 218100 696934
rect 222200 683188 222252 683194
rect 222200 683130 222252 683136
rect 222212 673454 222240 683130
rect 227168 676864 227220 676870
rect 227168 676806 227220 676812
rect 222212 673426 222424 673454
rect 222396 669882 222424 673426
rect 227180 669882 227208 676806
rect 232688 675504 232740 675510
rect 232688 675446 232740 675452
rect 232700 669882 232728 675446
rect 234632 674354 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 264980 700868 265032 700874
rect 264980 700810 265032 700816
rect 249800 700664 249852 700670
rect 249800 700606 249852 700612
rect 236000 700460 236052 700466
rect 236000 700402 236052 700408
rect 236012 692774 236040 700402
rect 249812 692774 249840 700606
rect 236012 692746 236592 692774
rect 249812 692746 250760 692774
rect 234620 674348 234672 674354
rect 234620 674290 234672 674296
rect 218072 669854 218178 669882
rect 222396 669854 222870 669882
rect 227180 669854 227562 669882
rect 232346 669854 232728 669882
rect 236564 669882 236592 692746
rect 241520 676932 241572 676938
rect 241520 676874 241572 676880
rect 241532 669882 241560 676874
rect 246672 675572 246724 675578
rect 246672 675514 246724 675520
rect 246684 669882 246712 675514
rect 236564 669854 237038 669882
rect 241532 669854 241730 669882
rect 246422 669854 246712 669882
rect 250732 669882 250760 692746
rect 255320 677000 255372 677006
rect 255320 676942 255372 676948
rect 255332 669882 255360 676942
rect 260656 675640 260708 675646
rect 260656 675582 260708 675588
rect 260668 669882 260696 675582
rect 250732 669854 251114 669882
rect 255332 669854 255806 669882
rect 260498 669854 260696 669882
rect 264992 669882 265020 700810
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 266372 675782 266400 697546
rect 282932 677278 282960 702406
rect 282920 677272 282972 677278
rect 282920 677214 282972 677220
rect 292856 677272 292908 677278
rect 292856 677214 292908 677220
rect 278872 677204 278924 677210
rect 278872 677146 278924 677152
rect 269488 677136 269540 677142
rect 269488 677078 269540 677084
rect 266360 675776 266412 675782
rect 266360 675718 266412 675724
rect 269500 669882 269528 677078
rect 274456 675708 274508 675714
rect 274456 675650 274508 675656
rect 274468 669882 274496 675650
rect 278884 669882 278912 677146
rect 288440 675776 288492 675782
rect 288440 675718 288492 675724
rect 284208 674416 284260 674422
rect 284208 674358 284260 674364
rect 284220 669882 284248 674358
rect 264992 669854 265190 669882
rect 269500 669854 269882 669882
rect 274468 669854 274574 669882
rect 278884 669854 279266 669882
rect 283958 669854 284248 669882
rect 288452 669882 288480 675718
rect 292868 669882 292896 677214
rect 299492 674422 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 306380 700936 306432 700942
rect 306380 700878 306432 700884
rect 306392 692774 306420 700878
rect 320180 700800 320232 700806
rect 320180 700742 320232 700748
rect 316040 700732 316092 700738
rect 316040 700674 316092 700680
rect 316052 692774 316080 700674
rect 320192 692774 320220 700742
rect 329840 700528 329892 700534
rect 329840 700470 329892 700476
rect 329852 692774 329880 700470
rect 306392 692746 307064 692774
rect 316052 692746 316448 692774
rect 320192 692746 321048 692774
rect 329852 692746 330432 692774
rect 302240 677068 302292 677074
rect 302240 677010 302292 677016
rect 299480 674416 299532 674422
rect 299480 674358 299532 674364
rect 297732 674348 297784 674354
rect 297732 674290 297784 674296
rect 297744 669882 297772 674290
rect 302252 669882 302280 677010
rect 307036 669882 307064 692746
rect 311900 674280 311952 674286
rect 311900 674222 311952 674228
rect 311912 669882 311940 674222
rect 316420 669882 316448 692746
rect 321020 669882 321048 692746
rect 325884 674212 325936 674218
rect 325884 674154 325936 674160
rect 325896 669882 325924 674154
rect 330404 669882 330432 692746
rect 331232 675714 331260 702986
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 335360 700596 335412 700602
rect 335360 700538 335412 700544
rect 331220 675708 331272 675714
rect 331220 675650 331272 675656
rect 335372 669882 335400 700538
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 345032 692774 345060 700266
rect 345032 692746 345152 692774
rect 340052 674144 340104 674150
rect 340052 674086 340104 674092
rect 340064 669882 340092 674086
rect 345124 669882 345152 692746
rect 347792 677210 347820 702406
rect 349160 700392 349212 700398
rect 349160 700334 349212 700340
rect 349172 692774 349200 700334
rect 349172 692746 349384 692774
rect 347780 677204 347832 677210
rect 347780 677146 347832 677152
rect 288452 669854 288650 669882
rect 292868 669854 293342 669882
rect 297744 669854 298034 669882
rect 302252 669854 302726 669882
rect 307036 669854 307418 669882
rect 311912 669854 312110 669882
rect 316420 669854 316802 669882
rect 321020 669854 321494 669882
rect 325896 669854 326186 669882
rect 330404 669854 330878 669882
rect 335372 669854 335570 669882
rect 340064 669854 340354 669882
rect 345046 669854 345152 669882
rect 349356 669882 349384 692746
rect 353944 683256 353996 683262
rect 353944 683198 353996 683204
rect 353956 669882 353984 683198
rect 364352 677142 364380 702406
rect 364340 677136 364392 677142
rect 364340 677078 364392 677084
rect 397472 675646 397500 703520
rect 413664 700874 413692 703520
rect 413652 700868 413704 700874
rect 413652 700810 413704 700816
rect 429212 677006 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 677000 429252 677006
rect 429200 676942 429252 676948
rect 397460 675640 397512 675646
rect 397460 675582 397512 675588
rect 462332 675578 462360 703520
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 494072 676938 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 676932 494112 676938
rect 494060 676874 494112 676880
rect 462320 675572 462372 675578
rect 462320 675514 462372 675520
rect 527192 675510 527220 703520
rect 543476 700466 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 558932 676870 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 558920 676864 558972 676870
rect 558920 676806 558972 676812
rect 527180 675504 527232 675510
rect 527180 675446 527232 675452
rect 557172 675436 557224 675442
rect 557172 675378 557224 675384
rect 556988 675368 557040 675374
rect 556988 675310 557040 675316
rect 555976 675300 556028 675306
rect 555976 675242 556028 675248
rect 555884 675232 555936 675238
rect 555884 675174 555936 675180
rect 555792 675164 555844 675170
rect 555792 675106 555844 675112
rect 554596 675096 554648 675102
rect 554596 675038 554648 675044
rect 554412 675028 554464 675034
rect 554412 674970 554464 674976
rect 513748 674892 513800 674898
rect 513748 674834 513800 674840
rect 368572 674008 368624 674014
rect 368572 673950 368624 673956
rect 363420 671492 363472 671498
rect 363420 671434 363472 671440
rect 363432 669882 363460 671434
rect 368584 669882 368612 673950
rect 372804 673940 372856 673946
rect 372804 673882 372856 673888
rect 349356 669854 349738 669882
rect 353956 669854 354430 669882
rect 363432 669854 363814 669882
rect 368506 669854 368612 669882
rect 372816 669882 372844 673882
rect 386972 673872 387024 673878
rect 386972 673814 387024 673820
rect 471426 673840 471482 673849
rect 377588 672988 377640 672994
rect 377588 672930 377640 672936
rect 377600 669882 377628 672930
rect 382280 671356 382332 671362
rect 382280 671298 382332 671304
rect 382292 669882 382320 671298
rect 386984 669882 387012 673814
rect 400956 673804 401008 673810
rect 471426 673775 471482 673784
rect 400956 673746 401008 673752
rect 392032 672920 392084 672926
rect 392032 672862 392084 672868
rect 395436 672920 395488 672926
rect 395436 672862 395488 672868
rect 392044 669882 392072 672862
rect 395448 670274 395476 672862
rect 397090 672480 397146 672489
rect 397090 672415 397146 672424
rect 397104 671362 397132 672415
rect 397092 671356 397144 671362
rect 397092 671298 397144 671304
rect 396354 671120 396410 671129
rect 396354 671055 396410 671064
rect 395436 670268 395488 670274
rect 395436 670210 395488 670216
rect 372816 669854 373198 669882
rect 377600 669854 377890 669882
rect 382292 669854 382582 669882
rect 386984 669854 387274 669882
rect 391966 669854 392072 669882
rect 396368 669882 396396 671055
rect 400968 669882 400996 673746
rect 415492 673736 415544 673742
rect 415492 673678 415544 673684
rect 405740 672852 405792 672858
rect 405740 672794 405792 672800
rect 405752 669882 405780 672794
rect 410340 671084 410392 671090
rect 410340 671026 410392 671032
rect 410352 669882 410380 671026
rect 415504 669882 415532 673678
rect 429200 673668 429252 673674
rect 429200 673610 429252 673616
rect 419724 672716 419776 672722
rect 419724 672658 419776 672664
rect 419816 672716 419868 672722
rect 419816 672658 419868 672664
rect 396368 669854 396658 669882
rect 400968 669854 401350 669882
rect 405752 669854 406042 669882
rect 410352 669854 410734 669882
rect 415426 669854 415532 669882
rect 419736 669882 419764 672658
rect 419828 670138 419856 672658
rect 424508 671016 424560 671022
rect 424508 670958 424560 670964
rect 419816 670132 419868 670138
rect 419816 670074 419868 670080
rect 424520 669882 424548 670958
rect 429212 669882 429240 673610
rect 443276 673600 443328 673606
rect 443276 673542 443328 673548
rect 433892 672580 433944 672586
rect 433892 672522 433944 672528
rect 433904 669882 433932 672522
rect 438950 670984 439006 670993
rect 438950 670919 439006 670928
rect 438964 669882 438992 670919
rect 419736 669854 420118 669882
rect 424520 669854 424810 669882
rect 429212 669854 429502 669882
rect 433904 669854 434194 669882
rect 438886 669854 438992 669882
rect 443288 669882 443316 673542
rect 457444 673532 457496 673538
rect 457444 673474 457496 673480
rect 452660 672920 452712 672926
rect 452660 672862 452712 672868
rect 448060 672444 448112 672450
rect 448060 672386 448112 672392
rect 448152 672444 448204 672450
rect 448152 672386 448204 672392
rect 448072 669882 448100 672386
rect 448164 670041 448192 672386
rect 448150 670032 448206 670041
rect 448150 669967 448206 669976
rect 452672 669882 452700 672862
rect 457456 669882 457484 673474
rect 462320 672376 462372 672382
rect 462320 672318 462372 672324
rect 462332 669882 462360 672318
rect 466828 670880 466880 670886
rect 466828 670822 466880 670828
rect 466840 669882 466868 670822
rect 471440 669882 471468 673775
rect 485778 673704 485834 673713
rect 485778 673639 485834 673648
rect 480812 672716 480864 672722
rect 480812 672658 480864 672664
rect 476212 672240 476264 672246
rect 476212 672182 476264 672188
rect 476224 669882 476252 672182
rect 480824 669882 480852 672658
rect 485792 669882 485820 673639
rect 499578 673568 499634 673577
rect 499578 673503 499634 673512
rect 490196 672172 490248 672178
rect 490196 672114 490248 672120
rect 490208 669882 490236 672114
rect 494980 670744 495032 670750
rect 494980 670686 495032 670692
rect 494992 669882 495020 670686
rect 499592 669882 499620 673503
rect 509240 672444 509292 672450
rect 509240 672386 509292 672392
rect 504364 672104 504416 672110
rect 504364 672046 504416 672052
rect 504376 669882 504404 672046
rect 509252 669882 509280 672386
rect 513760 669882 513788 674834
rect 532698 672616 532754 672625
rect 532698 672551 532754 672560
rect 518346 672344 518402 672353
rect 518346 672279 518402 672288
rect 518360 669882 518388 672279
rect 523130 671256 523186 671265
rect 523130 671191 523186 671200
rect 523144 669882 523172 671191
rect 532712 669882 532740 672551
rect 554136 672308 554188 672314
rect 554136 672250 554188 672256
rect 554044 670812 554096 670818
rect 554044 670754 554096 670760
rect 553952 670064 554004 670070
rect 553952 670006 554004 670012
rect 443288 669854 443578 669882
rect 448072 669854 448362 669882
rect 452672 669854 453054 669882
rect 457456 669854 457746 669882
rect 462332 669854 462438 669882
rect 466840 669854 467130 669882
rect 471440 669854 471822 669882
rect 476224 669854 476514 669882
rect 480824 669854 481206 669882
rect 485792 669854 485898 669882
rect 490208 669854 490590 669882
rect 494992 669854 495282 669882
rect 499592 669854 499974 669882
rect 504376 669854 504666 669882
rect 509252 669854 509358 669882
rect 513760 669854 514050 669882
rect 518360 669854 518742 669882
rect 523144 669854 523434 669882
rect 532712 669854 532818 669882
rect 139490 669624 139546 669633
rect 58558 669598 58860 669604
rect 58558 669582 58848 669598
rect 82018 669594 82400 669610
rect 82018 669588 82412 669594
rect 82018 669582 82360 669588
rect 162122 669624 162178 669633
rect 161874 669582 162122 669610
rect 139490 669559 139546 669568
rect 162122 669559 162178 669568
rect 358910 669624 358966 669633
rect 358966 669582 359122 669610
rect 358910 669559 358966 669568
rect 82360 669530 82412 669536
rect 77576 669520 77628 669526
rect 35438 669488 35494 669497
rect 35098 669446 35438 669474
rect 63250 669458 63448 669474
rect 77326 669468 77576 669474
rect 77326 669462 77628 669468
rect 63250 669452 63460 669458
rect 63250 669446 63408 669452
rect 35438 669423 35494 669432
rect 77326 669446 77616 669462
rect 63408 669394 63460 669400
rect 49424 669384 49476 669390
rect 16486 669352 16542 669361
rect 16330 669310 16486 669338
rect 21270 669352 21326 669361
rect 21022 669310 21270 669338
rect 16486 669287 16542 669296
rect 25962 669352 26018 669361
rect 25714 669310 25962 669338
rect 21270 669287 21326 669296
rect 30654 669352 30710 669361
rect 30406 669310 30654 669338
rect 25962 669287 26018 669296
rect 39946 669352 40002 669361
rect 39790 669310 39946 669338
rect 30654 669287 30710 669296
rect 49174 669332 49424 669338
rect 49174 669326 49476 669332
rect 527730 669352 527786 669361
rect 49174 669310 49464 669326
rect 39946 669287 40002 669296
rect 537114 669352 537170 669361
rect 527786 669310 528126 669338
rect 527730 669287 527786 669296
rect 541898 669352 541954 669361
rect 537170 669310 537510 669338
rect 537114 669287 537170 669296
rect 546590 669352 546646 669361
rect 541954 669310 542202 669338
rect 541898 669287 541954 669296
rect 546646 669310 546894 669338
rect 546590 669287 546646 669296
rect 13832 634786 13952 634814
rect 13832 633418 13860 634786
rect 13820 633412 13872 633418
rect 13820 633354 13872 633360
rect 553964 592006 553992 670006
rect 553952 592000 554004 592006
rect 553952 591942 554004 591948
rect 13360 580984 13412 580990
rect 13360 580926 13412 580932
rect 13268 476060 13320 476066
rect 13268 476002 13320 476008
rect 13176 423632 13228 423638
rect 13176 423574 13228 423580
rect 13084 411256 13136 411262
rect 13084 411198 13136 411204
rect 554056 167006 554084 670754
rect 554148 219434 554176 672250
rect 554228 669860 554280 669866
rect 554228 669802 554280 669808
rect 554240 259418 554268 669802
rect 554320 669792 554372 669798
rect 554320 669734 554372 669740
rect 554332 273222 554360 669734
rect 554424 325650 554452 674970
rect 554504 670948 554556 670954
rect 554504 670890 554556 670896
rect 554516 353258 554544 670890
rect 554608 379506 554636 675038
rect 555700 672784 555752 672790
rect 555700 672726 555752 672732
rect 555608 672648 555660 672654
rect 555608 672590 555660 672596
rect 555516 672512 555568 672518
rect 555516 672454 555568 672460
rect 555332 670200 555384 670206
rect 555332 670142 555384 670148
rect 554688 669928 554740 669934
rect 554688 669870 554740 669876
rect 554700 405686 554728 669870
rect 555344 632058 555372 670142
rect 555424 669656 555476 669662
rect 555424 669598 555476 669604
rect 555332 632052 555384 632058
rect 555332 631994 555384 632000
rect 554688 405680 554740 405686
rect 554688 405622 554740 405628
rect 554596 379500 554648 379506
rect 554596 379442 554648 379448
rect 554504 353252 554556 353258
rect 554504 353194 554556 353200
rect 554412 325644 554464 325650
rect 554412 325586 554464 325592
rect 554320 273216 554372 273222
rect 554320 273158 554372 273164
rect 554228 259412 554280 259418
rect 554228 259354 554280 259360
rect 554136 219428 554188 219434
rect 554136 219370 554188 219376
rect 554044 167000 554096 167006
rect 554044 166942 554096 166948
rect 11704 137964 11756 137970
rect 11704 137906 11756 137912
rect 555436 126954 555464 669598
rect 555528 313274 555556 672454
rect 555620 365702 555648 672590
rect 555712 419490 555740 672726
rect 555804 431934 555832 675106
rect 555896 458182 555924 675174
rect 555988 471986 556016 675242
rect 556802 673976 556858 673985
rect 556802 673911 556858 673920
rect 556068 671288 556120 671294
rect 556068 671230 556120 671236
rect 556080 564398 556108 671230
rect 556068 564392 556120 564398
rect 556068 564334 556120 564340
rect 555976 471980 556028 471986
rect 555976 471922 556028 471928
rect 555884 458176 555936 458182
rect 555884 458118 555936 458124
rect 555792 431928 555844 431934
rect 555792 431870 555844 431876
rect 555700 419484 555752 419490
rect 555700 419426 555752 419432
rect 555608 365696 555660 365702
rect 555608 365638 555660 365644
rect 555516 313268 555568 313274
rect 555516 313210 555568 313216
rect 556816 245614 556844 673911
rect 556896 671152 556948 671158
rect 556896 671094 556948 671100
rect 556908 511970 556936 671094
rect 557000 525774 557028 675310
rect 557080 671220 557132 671226
rect 557080 671162 557132 671168
rect 557092 538218 557120 671162
rect 557184 578202 557212 675378
rect 580172 674960 580224 674966
rect 580172 674902 580224 674908
rect 557356 674076 557408 674082
rect 557356 674018 557408 674024
rect 557264 671560 557316 671566
rect 557264 671502 557316 671508
rect 557276 618254 557304 671502
rect 557368 644434 557396 674018
rect 579620 671424 579672 671430
rect 579620 671366 579672 671372
rect 579632 670721 579660 671366
rect 579618 670712 579674 670721
rect 579618 670647 579674 670656
rect 580078 668536 580134 668545
rect 580078 668471 580134 668480
rect 557356 644428 557408 644434
rect 557356 644370 557408 644376
rect 579988 644428 580040 644434
rect 579988 644370 580040 644376
rect 580000 644065 580028 644370
rect 579986 644056 580042 644065
rect 579986 643991 580042 644000
rect 579988 632052 580040 632058
rect 579988 631994 580040 632000
rect 580000 630873 580028 631994
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 557264 618248 557316 618254
rect 557264 618190 557316 618196
rect 579988 618248 580040 618254
rect 579988 618190 580040 618196
rect 580000 617545 580028 618190
rect 579986 617536 580042 617545
rect 579986 617471 580042 617480
rect 579804 592000 579856 592006
rect 579804 591942 579856 591948
rect 579816 591025 579844 591942
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 557172 578196 557224 578202
rect 557172 578138 557224 578144
rect 579804 578196 579856 578202
rect 579804 578138 579856 578144
rect 579816 577697 579844 578138
rect 579802 577688 579858 577697
rect 579802 577623 579858 577632
rect 579988 564392 580040 564398
rect 579986 564360 579988 564369
rect 580040 564360 580042 564369
rect 579986 564295 580042 564304
rect 557080 538212 557132 538218
rect 557080 538154 557132 538160
rect 579988 538212 580040 538218
rect 579988 538154 580040 538160
rect 580000 537849 580028 538154
rect 579986 537840 580042 537849
rect 579986 537775 580042 537784
rect 556988 525768 557040 525774
rect 556988 525710 557040 525716
rect 579988 525768 580040 525774
rect 579988 525710 580040 525716
rect 580000 524521 580028 525710
rect 579986 524512 580042 524521
rect 579986 524447 580042 524456
rect 556896 511964 556948 511970
rect 556896 511906 556948 511912
rect 579988 511964 580040 511970
rect 579988 511906 580040 511912
rect 580000 511329 580028 511906
rect 579986 511320 580042 511329
rect 579986 511255 580042 511264
rect 579804 471980 579856 471986
rect 579804 471922 579856 471928
rect 579816 471481 579844 471922
rect 579802 471472 579858 471481
rect 579802 471407 579858 471416
rect 579988 458176 580040 458182
rect 579986 458144 579988 458153
rect 580040 458144 580042 458153
rect 579986 458079 580042 458088
rect 579988 431928 580040 431934
rect 579988 431870 580040 431876
rect 580000 431633 580028 431870
rect 579986 431624 580042 431633
rect 579986 431559 580042 431568
rect 579988 419484 580040 419490
rect 579988 419426 580040 419432
rect 580000 418305 580028 419426
rect 579986 418296 580042 418305
rect 579986 418231 580042 418240
rect 579988 405680 580040 405686
rect 579988 405622 580040 405628
rect 580000 404977 580028 405622
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 579804 379500 579856 379506
rect 579804 379442 579856 379448
rect 579816 378457 579844 379442
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579988 365696 580040 365702
rect 579988 365638 580040 365644
rect 580000 365129 580028 365638
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 579988 353252 580040 353258
rect 579988 353194 580040 353200
rect 580000 351937 580028 353194
rect 579986 351928 580042 351937
rect 579986 351863 580042 351872
rect 579988 325644 580040 325650
rect 579988 325586 580040 325592
rect 580000 325281 580028 325586
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 579988 313268 580040 313274
rect 579988 313210 580040 313216
rect 580000 312089 580028 313210
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580092 298761 580120 668471
rect 580078 298752 580134 298761
rect 580078 298687 580134 298696
rect 580080 273216 580132 273222
rect 580080 273158 580132 273164
rect 580092 272241 580120 273158
rect 580078 272232 580134 272241
rect 580078 272167 580134 272176
rect 580080 259412 580132 259418
rect 580080 259354 580132 259360
rect 580092 258913 580120 259354
rect 580078 258904 580134 258913
rect 580078 258839 580134 258848
rect 556804 245608 556856 245614
rect 580080 245608 580132 245614
rect 556804 245550 556856 245556
rect 580078 245576 580080 245585
rect 580132 245576 580134 245585
rect 580078 245511 580134 245520
rect 580184 232393 580212 674902
rect 580540 671356 580592 671362
rect 580540 671298 580592 671304
rect 580356 669996 580408 670002
rect 580356 669938 580408 669944
rect 580262 669352 580318 669361
rect 580262 669287 580318 669296
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579620 167000 579672 167006
rect 579620 166942 579672 166948
rect 579632 165889 579660 166942
rect 579618 165880 579674 165889
rect 579618 165815 579674 165824
rect 555424 126948 555476 126954
rect 555424 126890 555476 126896
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 4988 97912 5040 97918
rect 4988 97854 5040 97860
rect 4896 84924 4948 84930
rect 4896 84866 4948 84872
rect 580276 59673 580304 669287
rect 580368 99521 580396 669938
rect 580448 669384 580500 669390
rect 580448 669326 580500 669332
rect 580460 112849 580488 669326
rect 580552 139369 580580 671298
rect 580908 669724 580960 669730
rect 580908 669666 580960 669672
rect 580724 669588 580776 669594
rect 580724 669530 580776 669536
rect 580632 669452 580684 669458
rect 580632 669394 580684 669400
rect 580644 152697 580672 669394
rect 580736 179217 580764 669530
rect 580816 669520 580868 669526
rect 580816 669462 580868 669468
rect 580828 192545 580856 669462
rect 580920 205737 580948 669666
rect 580906 205728 580962 205737
rect 580906 205663 580962 205672
rect 580814 192536 580870 192545
rect 580814 192471 580870 192480
rect 580722 179208 580778 179217
rect 580722 179143 580778 179152
rect 580630 152688 580686 152697
rect 580630 152623 580686 152632
rect 580538 139360 580594 139369
rect 580538 139295 580594 139304
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580354 99512 580410 99521
rect 580354 99447 580410 99456
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 2780 58676 2832 58682
rect 2780 58618 2832 58624
rect 4804 58676 4856 58682
rect 4804 58618 4856 58624
rect 2792 58585 2820 58618
rect 2778 58576 2834 58585
rect 2778 58511 2834 58520
rect 13832 50102 14490 50130
rect 15304 50102 15502 50130
rect 16606 50102 16712 50130
rect 11060 48204 11112 48210
rect 11060 48146 11112 48152
rect 2780 47864 2832 47870
rect 2780 47806 2832 47812
rect 2792 16574 2820 47806
rect 8300 47796 8352 47802
rect 8300 47738 8352 47744
rect 6920 47728 6972 47734
rect 6920 47670 6972 47676
rect 5540 47660 5592 47666
rect 5540 47602 5592 47608
rect 4160 47592 4212 47598
rect 4160 47534 4212 47540
rect 4172 16574 4200 47534
rect 5552 16574 5580 47602
rect 6932 16574 6960 47670
rect 8312 16574 8340 47738
rect 9680 47524 9732 47530
rect 9680 47466 9732 47472
rect 2792 16546 3648 16574
rect 4172 16546 5304 16574
rect 5552 16546 6040 16574
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 47466
rect 11072 6914 11100 48146
rect 11152 48000 11204 48006
rect 11152 47942 11204 47948
rect 11164 16574 11192 47942
rect 12440 47932 12492 47938
rect 12440 47874 12492 47880
rect 12452 16574 12480 47874
rect 11164 16546 11928 16574
rect 12452 16546 13584 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13556 480 13584 16546
rect 13832 3466 13860 50102
rect 15200 48068 15252 48074
rect 15200 48010 15252 48016
rect 13912 47388 13964 47394
rect 13912 47330 13964 47336
rect 13924 16574 13952 47330
rect 13924 16546 14320 16574
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15212 3482 15240 48010
rect 15304 3602 15332 50102
rect 16580 48136 16632 48142
rect 16580 48078 16632 48084
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 16592 3482 16620 48078
rect 16684 3602 16712 50102
rect 17328 50102 17710 50130
rect 18432 50102 18814 50130
rect 19536 50102 19918 50130
rect 20732 50102 21022 50130
rect 22126 50102 22232 50130
rect 17328 47870 17356 50102
rect 17316 47864 17368 47870
rect 17316 47806 17368 47812
rect 18432 47598 18460 50102
rect 19536 47666 19564 50102
rect 19616 47864 19668 47870
rect 19616 47806 19668 47812
rect 19524 47660 19576 47666
rect 19524 47602 19576 47608
rect 18420 47592 18472 47598
rect 18420 47534 18472 47540
rect 17960 47456 18012 47462
rect 17960 47398 18012 47404
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 15212 3454 15976 3482
rect 16592 3454 17080 3482
rect 15948 480 15976 3454
rect 17052 480 17080 3454
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 47398
rect 19628 45554 19656 47806
rect 20732 47734 20760 50102
rect 22204 47802 22232 50102
rect 22848 50102 23230 50130
rect 23952 50102 24334 50130
rect 25056 50102 25438 50130
rect 26344 50102 26450 50130
rect 27264 50102 27554 50130
rect 28368 50102 28658 50130
rect 29472 50102 29762 50130
rect 30576 50102 30866 50130
rect 31772 50102 31970 50130
rect 32784 50102 33074 50130
rect 33888 50102 34178 50130
rect 34992 50102 35282 50130
rect 36096 50102 36386 50130
rect 37292 50102 37490 50130
rect 38120 50102 38502 50130
rect 39224 50102 39606 50130
rect 40328 50102 40710 50130
rect 41432 50102 41814 50130
rect 42918 50102 43024 50130
rect 22284 48272 22336 48278
rect 22284 48214 22336 48220
rect 22192 47796 22244 47802
rect 22192 47738 22244 47744
rect 20720 47728 20772 47734
rect 20720 47670 20772 47676
rect 20720 47592 20772 47598
rect 20720 47534 20772 47540
rect 19536 45526 19656 45554
rect 19536 6914 19564 45526
rect 20732 16574 20760 47534
rect 22296 16574 22324 48214
rect 22848 47530 22876 50102
rect 23952 48210 23980 50102
rect 23940 48204 23992 48210
rect 23940 48146 23992 48152
rect 24952 48204 25004 48210
rect 24952 48146 25004 48152
rect 23480 47796 23532 47802
rect 23480 47738 23532 47744
rect 22836 47524 22888 47530
rect 22836 47466 22888 47472
rect 23492 16574 23520 47738
rect 24964 16574 24992 48146
rect 25056 48006 25084 50102
rect 25044 48000 25096 48006
rect 25044 47942 25096 47948
rect 26344 47938 26372 50102
rect 26332 47932 26384 47938
rect 26332 47874 26384 47880
rect 26240 47524 26292 47530
rect 26240 47466 26292 47472
rect 25504 47252 25556 47258
rect 25504 47194 25556 47200
rect 20732 16546 21864 16574
rect 22296 16546 22600 16574
rect 23492 16546 24256 16574
rect 24964 16546 25360 16574
rect 19444 6886 19564 6914
rect 19444 480 19472 6886
rect 20628 3324 20680 3330
rect 20628 3266 20680 3272
rect 20640 480 20668 3266
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 25516 3330 25544 47194
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 47466
rect 27264 47394 27292 50102
rect 28368 48074 28396 50102
rect 29472 48142 29500 50102
rect 29460 48136 29512 48142
rect 29460 48078 29512 48084
rect 28356 48068 28408 48074
rect 28356 48010 28408 48016
rect 27620 47728 27672 47734
rect 27620 47670 27672 47676
rect 27252 47388 27304 47394
rect 27252 47330 27304 47336
rect 27632 3534 27660 47670
rect 29000 47660 29052 47666
rect 29000 47602 29052 47608
rect 27712 47320 27764 47326
rect 27712 47262 27764 47268
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27724 480 27752 47262
rect 29012 16574 29040 47602
rect 30576 47462 30604 50102
rect 31772 47870 31800 50102
rect 31944 48000 31996 48006
rect 31944 47942 31996 47948
rect 31760 47864 31812 47870
rect 31760 47806 31812 47812
rect 30564 47456 30616 47462
rect 30564 47398 30616 47404
rect 29012 16546 30144 16574
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3470
rect 30116 480 30144 16546
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31312 480 31340 3402
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 47942
rect 32784 47258 32812 50102
rect 33232 47932 33284 47938
rect 33232 47874 33284 47880
rect 32772 47252 32824 47258
rect 32772 47194 32824 47200
rect 33244 16574 33272 47874
rect 33888 47598 33916 50102
rect 34992 48278 35020 50102
rect 34980 48272 35032 48278
rect 34980 48214 35032 48220
rect 35992 48272 36044 48278
rect 35992 48214 36044 48220
rect 33876 47592 33928 47598
rect 33876 47534 33928 47540
rect 35900 47592 35952 47598
rect 35900 47534 35952 47540
rect 34520 47456 34572 47462
rect 34520 47398 34572 47404
rect 33244 16546 33640 16574
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 47398
rect 35912 3534 35940 47534
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 48214
rect 36096 47802 36124 50102
rect 37292 48210 37320 50102
rect 37280 48204 37332 48210
rect 37280 48146 37332 48152
rect 36084 47796 36136 47802
rect 36084 47738 36136 47744
rect 38120 47530 38148 50102
rect 38752 48068 38804 48074
rect 38752 48010 38804 48016
rect 38108 47524 38160 47530
rect 38108 47466 38160 47472
rect 37280 47388 37332 47394
rect 37280 47330 37332 47336
rect 37292 16574 37320 47330
rect 38764 16574 38792 48010
rect 39224 47326 39252 50102
rect 40132 47864 40184 47870
rect 40132 47806 40184 47812
rect 39212 47320 39264 47326
rect 39212 47262 39264 47268
rect 40144 16574 40172 47806
rect 40328 47734 40356 50102
rect 40316 47728 40368 47734
rect 40316 47670 40368 47676
rect 41432 47666 41460 50102
rect 41512 48204 41564 48210
rect 41512 48146 41564 48152
rect 41420 47660 41472 47666
rect 41420 47602 41472 47608
rect 41524 16574 41552 48146
rect 42800 47660 42852 47666
rect 42800 47602 42852 47608
rect 37292 16546 38424 16574
rect 38764 16546 39160 16574
rect 40144 16546 40264 16574
rect 41524 16546 41920 16574
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 47602
rect 42996 45554 43024 50102
rect 43640 50102 44022 50130
rect 44744 50102 45126 50130
rect 45848 50102 46230 50130
rect 46952 50102 47334 50130
rect 48332 50102 48438 50130
rect 49160 50102 49542 50130
rect 50264 50102 50554 50130
rect 51368 50102 51658 50130
rect 52472 50102 52762 50130
rect 53866 50102 53972 50130
rect 43640 48006 43668 50102
rect 44364 48136 44416 48142
rect 44364 48078 44416 48084
rect 43628 48000 43680 48006
rect 43628 47942 43680 47948
rect 44272 47320 44324 47326
rect 44272 47262 44324 47268
rect 42904 45526 43024 45554
rect 42904 3466 42932 45526
rect 42892 3460 42944 3466
rect 42892 3402 42944 3408
rect 44284 480 44312 47262
rect 44376 16574 44404 48078
rect 44744 47938 44772 50102
rect 44732 47932 44784 47938
rect 44732 47874 44784 47880
rect 45652 47932 45704 47938
rect 45652 47874 45704 47880
rect 45664 16574 45692 47874
rect 45848 47462 45876 50102
rect 46952 48278 46980 50102
rect 46940 48272 46992 48278
rect 46940 48214 46992 48220
rect 46940 47796 46992 47802
rect 46940 47738 46992 47744
rect 45836 47456 45888 47462
rect 45836 47398 45888 47404
rect 46952 16574 46980 47738
rect 48332 47598 48360 50102
rect 48412 47728 48464 47734
rect 48412 47670 48464 47676
rect 48320 47592 48372 47598
rect 48320 47534 48372 47540
rect 48424 16574 48452 47670
rect 49160 47394 49188 50102
rect 50264 48074 50292 50102
rect 50252 48068 50304 48074
rect 50252 48010 50304 48016
rect 51172 48000 51224 48006
rect 51172 47942 51224 47948
rect 49700 47524 49752 47530
rect 49700 47466 49752 47472
rect 49148 47388 49200 47394
rect 49148 47330 49200 47336
rect 49712 16574 49740 47466
rect 44376 16546 45048 16574
rect 45664 16546 46704 16574
rect 46952 16546 47440 16574
rect 48424 16546 48544 16574
rect 49712 16546 50200 16574
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51184 354 51212 47942
rect 51368 47870 51396 50102
rect 52472 48210 52500 50102
rect 52460 48204 52512 48210
rect 52460 48146 52512 48152
rect 52552 48204 52604 48210
rect 52552 48146 52604 48152
rect 51356 47864 51408 47870
rect 51356 47806 51408 47812
rect 52460 47592 52512 47598
rect 52460 47534 52512 47540
rect 52472 3534 52500 47534
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 48146
rect 53944 47666 53972 50102
rect 54680 50102 54970 50130
rect 55784 50102 56074 50130
rect 56888 50102 57178 50130
rect 57992 50102 58282 50130
rect 59386 50102 59492 50130
rect 54024 47864 54076 47870
rect 54024 47806 54076 47812
rect 53932 47660 53984 47666
rect 53932 47602 53984 47608
rect 54036 16574 54064 47806
rect 54680 47326 54708 50102
rect 55312 48272 55364 48278
rect 55312 48214 55364 48220
rect 54668 47320 54720 47326
rect 54668 47262 54720 47268
rect 55324 16574 55352 48214
rect 55784 48142 55812 50102
rect 55772 48136 55824 48142
rect 55772 48078 55824 48084
rect 56692 48068 56744 48074
rect 56692 48010 56744 48016
rect 56704 16574 56732 48010
rect 56888 47938 56916 50102
rect 56876 47932 56928 47938
rect 56876 47874 56928 47880
rect 57992 47802 58020 50102
rect 57980 47796 58032 47802
rect 57980 47738 58032 47744
rect 59464 47734 59492 50102
rect 60200 50102 60490 50130
rect 61120 50102 61502 50130
rect 62224 50102 62606 50130
rect 63512 50102 63710 50130
rect 64432 50102 64814 50130
rect 65536 50102 65918 50130
rect 66640 50102 67022 50130
rect 67744 50102 68126 50130
rect 69032 50102 69230 50130
rect 69952 50102 70334 50130
rect 71056 50102 71438 50130
rect 72160 50102 72542 50130
rect 73264 50102 73554 50130
rect 74552 50102 74658 50130
rect 75472 50102 75762 50130
rect 76576 50102 76866 50130
rect 77680 50102 77970 50130
rect 78876 50102 79074 50130
rect 80072 50102 80178 50130
rect 80992 50102 81282 50130
rect 82096 50102 82386 50130
rect 83200 50102 83490 50130
rect 84304 50102 84594 50130
rect 85606 50102 85712 50130
rect 59544 47932 59596 47938
rect 59544 47874 59596 47880
rect 59452 47728 59504 47734
rect 59452 47670 59504 47676
rect 57980 47660 58032 47666
rect 57980 47602 58032 47608
rect 57992 16574 58020 47602
rect 59556 16574 59584 47874
rect 60200 47530 60228 50102
rect 60832 48136 60884 48142
rect 60832 48078 60884 48084
rect 60740 47796 60792 47802
rect 60740 47738 60792 47744
rect 60188 47524 60240 47530
rect 60188 47466 60240 47472
rect 54036 16546 54984 16574
rect 55324 16546 56088 16574
rect 56704 16546 56824 16574
rect 57992 16546 58480 16574
rect 59556 16546 59676 16574
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 51326 354 51438 480
rect 51184 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 59648 480 59676 16546
rect 60752 6914 60780 47738
rect 60844 16574 60872 48078
rect 61120 48006 61148 50102
rect 62224 48210 62252 50102
rect 62212 48204 62264 48210
rect 62212 48146 62264 48152
rect 61108 48000 61160 48006
rect 61108 47942 61160 47948
rect 62120 47728 62172 47734
rect 62120 47670 62172 47676
rect 62132 16574 62160 47670
rect 63512 47598 63540 50102
rect 63684 48000 63736 48006
rect 63684 47942 63736 47948
rect 63500 47592 63552 47598
rect 63500 47534 63552 47540
rect 63696 16574 63724 47942
rect 64432 47870 64460 50102
rect 65536 48278 65564 50102
rect 65524 48272 65576 48278
rect 65524 48214 65576 48220
rect 66640 48074 66668 50102
rect 66628 48068 66680 48074
rect 66628 48010 66680 48016
rect 64420 47864 64472 47870
rect 64420 47806 64472 47812
rect 67744 47666 67772 50102
rect 68284 48272 68336 48278
rect 68284 48214 68336 48220
rect 67824 47864 67876 47870
rect 67824 47806 67876 47812
rect 67732 47660 67784 47666
rect 67732 47602 67784 47608
rect 64880 47592 64932 47598
rect 64880 47534 64932 47540
rect 64892 16574 64920 47534
rect 67836 45554 67864 47806
rect 67744 45526 67864 45554
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 63696 16546 64368 16574
rect 64892 16546 65104 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 66732 480 66760 3470
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67744 354 67772 45526
rect 68296 3534 68324 48214
rect 69032 47938 69060 50102
rect 69112 48068 69164 48074
rect 69112 48010 69164 48016
rect 69020 47932 69072 47938
rect 69020 47874 69072 47880
rect 69020 47660 69072 47666
rect 69020 47602 69072 47608
rect 69032 3534 69060 47602
rect 68284 3528 68336 3534
rect 68284 3470 68336 3476
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 69124 480 69152 48010
rect 69952 47802 69980 50102
rect 71056 48142 71084 50102
rect 71044 48136 71096 48142
rect 71044 48078 71096 48084
rect 71872 47932 71924 47938
rect 71872 47874 71924 47880
rect 69940 47796 69992 47802
rect 69940 47738 69992 47744
rect 70400 47796 70452 47802
rect 70400 47738 70452 47744
rect 70412 16574 70440 47738
rect 71884 16574 71912 47874
rect 72160 47734 72188 50102
rect 73264 48006 73292 50102
rect 73252 48000 73304 48006
rect 73252 47942 73304 47948
rect 72148 47728 72200 47734
rect 72148 47670 72200 47676
rect 74552 47598 74580 50102
rect 75472 48278 75500 50102
rect 75460 48272 75512 48278
rect 75460 48214 75512 48220
rect 76576 47870 76604 50102
rect 77680 48074 77708 50102
rect 77668 48068 77720 48074
rect 77668 48010 77720 48016
rect 78772 48000 78824 48006
rect 78772 47942 78824 47948
rect 76564 47864 76616 47870
rect 76564 47806 76616 47812
rect 75920 47728 75972 47734
rect 75920 47670 75972 47676
rect 74540 47592 74592 47598
rect 74540 47534 74592 47540
rect 75184 47592 75236 47598
rect 75184 47534 75236 47540
rect 74540 47456 74592 47462
rect 74540 47398 74592 47404
rect 74552 16574 74580 47398
rect 70412 16546 71544 16574
rect 71884 16546 72648 16574
rect 74552 16546 75040 16574
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 67886 354 67998 480
rect 67744 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3470
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 73804 2984 73856 2990
rect 73804 2926 73856 2932
rect 73816 480 73844 2926
rect 75012 480 75040 16546
rect 75196 2990 75224 47534
rect 75184 2984 75236 2990
rect 75184 2926 75236 2932
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 47670
rect 77300 46980 77352 46986
rect 77300 46922 77352 46928
rect 77312 16574 77340 46922
rect 78784 16574 78812 47942
rect 78876 47666 78904 50102
rect 80072 47802 80100 50102
rect 80244 48068 80296 48074
rect 80244 48010 80296 48016
rect 80060 47796 80112 47802
rect 80060 47738 80112 47744
rect 78864 47660 78916 47666
rect 78864 47602 78916 47608
rect 80256 16574 80284 48010
rect 80992 47938 81020 50102
rect 80980 47932 81032 47938
rect 80980 47874 81032 47880
rect 81440 47660 81492 47666
rect 81440 47602 81492 47608
rect 81452 16574 81480 47602
rect 82096 47598 82124 50102
rect 82084 47592 82136 47598
rect 82084 47534 82136 47540
rect 82820 47592 82872 47598
rect 82820 47534 82872 47540
rect 82832 16574 82860 47534
rect 83200 47462 83228 50102
rect 84304 47734 84332 50102
rect 84292 47728 84344 47734
rect 84292 47670 84344 47676
rect 84292 47524 84344 47530
rect 84292 47466 84344 47472
rect 83188 47456 83240 47462
rect 83188 47398 83240 47404
rect 77312 16546 78168 16574
rect 78784 16546 79272 16574
rect 80256 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77392 4140 77444 4146
rect 77392 4082 77444 4088
rect 77404 480 77432 4082
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84304 354 84332 47466
rect 85580 47320 85632 47326
rect 85580 47262 85632 47268
rect 85592 6914 85620 47262
rect 85684 11778 85712 50102
rect 86328 50102 86710 50130
rect 87432 50102 87814 50130
rect 88536 50102 88918 50130
rect 89732 50102 90022 50130
rect 91126 50102 91232 50130
rect 85764 47864 85816 47870
rect 85764 47806 85816 47812
rect 85776 16574 85804 47806
rect 86328 46986 86356 50102
rect 87432 48006 87460 50102
rect 88536 48074 88564 50102
rect 88524 48068 88576 48074
rect 88524 48010 88576 48016
rect 87420 48000 87472 48006
rect 87420 47942 87472 47948
rect 86960 47796 87012 47802
rect 86960 47738 87012 47744
rect 86316 46980 86368 46986
rect 86316 46922 86368 46928
rect 86972 16574 87000 47738
rect 88340 47728 88392 47734
rect 88340 47670 88392 47676
rect 88352 16574 88380 47670
rect 89732 47666 89760 50102
rect 91100 48068 91152 48074
rect 91100 48010 91152 48016
rect 89812 48000 89864 48006
rect 89812 47942 89864 47948
rect 89720 47660 89772 47666
rect 89720 47602 89772 47608
rect 89824 16574 89852 47942
rect 91112 16574 91140 48010
rect 91204 47598 91232 50102
rect 91848 50102 92230 50130
rect 92952 50102 93334 50130
rect 94056 50102 94438 50130
rect 95252 50102 95542 50130
rect 96646 50102 96752 50130
rect 91192 47592 91244 47598
rect 91192 47534 91244 47540
rect 91848 47530 91876 50102
rect 92480 47932 92532 47938
rect 92480 47874 92532 47880
rect 91836 47524 91888 47530
rect 91836 47466 91888 47472
rect 85776 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89824 16546 89944 16574
rect 91112 16546 91600 16574
rect 85684 11750 85804 11778
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 85776 4146 85804 11750
rect 85764 4140 85816 4146
rect 85764 4082 85816 4088
rect 84446 354 84558 480
rect 84304 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 47874
rect 92952 47326 92980 50102
rect 94056 47870 94084 50102
rect 94044 47864 94096 47870
rect 94044 47806 94096 47812
rect 95252 47802 95280 50102
rect 96620 48204 96672 48210
rect 96620 48146 96672 48152
rect 95240 47796 95292 47802
rect 95240 47738 95292 47744
rect 95240 47660 95292 47666
rect 95240 47602 95292 47608
rect 93952 47592 94004 47598
rect 93952 47534 94004 47540
rect 92940 47320 92992 47326
rect 92940 47262 92992 47268
rect 93860 47320 93912 47326
rect 93860 47262 93912 47268
rect 93872 6914 93900 47262
rect 93964 16574 93992 47534
rect 95252 16574 95280 47602
rect 96632 16574 96660 48146
rect 96724 47734 96752 50102
rect 97368 50102 97658 50130
rect 98472 50102 98762 50130
rect 99576 50102 99866 50130
rect 100772 50102 100970 50130
rect 101784 50102 102074 50130
rect 102888 50102 103178 50130
rect 103992 50102 104282 50130
rect 105096 50102 105386 50130
rect 106292 50102 106490 50130
rect 107304 50102 107594 50130
rect 108224 50102 108606 50130
rect 109328 50102 109710 50130
rect 110432 50102 110814 50130
rect 111812 50102 111918 50130
rect 112640 50102 113022 50130
rect 113744 50102 114126 50130
rect 114848 50102 115230 50130
rect 115952 50102 116334 50130
rect 117332 50102 117438 50130
rect 118160 50102 118542 50130
rect 119264 50102 119646 50130
rect 120368 50102 120658 50130
rect 121564 50102 121762 50130
rect 122866 50102 122972 50130
rect 97368 48006 97396 50102
rect 98472 48074 98500 50102
rect 98460 48068 98512 48074
rect 98460 48010 98512 48016
rect 97356 48000 97408 48006
rect 97356 47942 97408 47948
rect 99576 47938 99604 50102
rect 99564 47932 99616 47938
rect 99564 47874 99616 47880
rect 98092 47864 98144 47870
rect 98092 47806 98144 47812
rect 96712 47728 96764 47734
rect 96712 47670 96764 47676
rect 98104 16574 98132 47806
rect 99380 47796 99432 47802
rect 99380 47738 99432 47744
rect 99392 16574 99420 47738
rect 100772 47326 100800 50102
rect 100944 48272 100996 48278
rect 100944 48214 100996 48220
rect 100760 47320 100812 47326
rect 100760 47262 100812 47268
rect 100956 16574 100984 48214
rect 101784 47598 101812 50102
rect 102324 47728 102376 47734
rect 102324 47670 102376 47676
rect 101772 47592 101824 47598
rect 101772 47534 101824 47540
rect 102336 16574 102364 47670
rect 102888 47666 102916 50102
rect 103992 48210 104020 50102
rect 103980 48204 104032 48210
rect 103980 48146 104032 48152
rect 103520 48068 103572 48074
rect 103520 48010 103572 48016
rect 102876 47660 102928 47666
rect 102876 47602 102928 47608
rect 103532 16574 103560 48010
rect 104900 48000 104952 48006
rect 104900 47942 104952 47948
rect 104912 16574 104940 47942
rect 105096 47870 105124 50102
rect 105084 47864 105136 47870
rect 105084 47806 105136 47812
rect 105544 47864 105596 47870
rect 105544 47806 105596 47812
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98104 16546 98224 16574
rect 99392 16546 99880 16574
rect 100956 16546 101076 16574
rect 102336 16546 103376 16574
rect 103532 16546 104112 16574
rect 104912 16546 105492 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 101048 480 101076 16546
rect 102232 3868 102284 3874
rect 102232 3810 102284 3816
rect 102244 480 102272 3810
rect 103348 480 103376 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105464 3482 105492 16546
rect 105556 3874 105584 47806
rect 106292 47802 106320 50102
rect 107304 48278 107332 50102
rect 107292 48272 107344 48278
rect 107292 48214 107344 48220
rect 108224 47870 108252 50102
rect 109132 47932 109184 47938
rect 109132 47874 109184 47880
rect 108212 47864 108264 47870
rect 108212 47806 108264 47812
rect 106280 47796 106332 47802
rect 106280 47738 106332 47744
rect 107660 47796 107712 47802
rect 107660 47738 107712 47744
rect 106280 47660 106332 47666
rect 106280 47602 106332 47608
rect 106292 16574 106320 47602
rect 107672 16574 107700 47738
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 105544 3868 105596 3874
rect 105544 3810 105596 3816
rect 105464 3454 105768 3482
rect 105740 480 105768 3454
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109144 354 109172 47874
rect 109328 47734 109356 50102
rect 110432 48074 110460 50102
rect 110420 48068 110472 48074
rect 110420 48010 110472 48016
rect 111812 48006 111840 50102
rect 111984 48068 112036 48074
rect 111984 48010 112036 48016
rect 111800 48000 111852 48006
rect 111800 47942 111852 47948
rect 109316 47728 109368 47734
rect 109316 47670 109368 47676
rect 110604 47728 110656 47734
rect 110604 47670 110656 47676
rect 110512 47592 110564 47598
rect 110512 47534 110564 47540
rect 110524 3534 110552 47534
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 110616 3346 110644 47670
rect 111996 16574 112024 48010
rect 112640 47666 112668 50102
rect 113180 48000 113232 48006
rect 113180 47942 113232 47948
rect 112628 47660 112680 47666
rect 112628 47602 112680 47608
rect 113192 16574 113220 47942
rect 113744 47802 113772 50102
rect 114848 47938 114876 50102
rect 114836 47932 114888 47938
rect 114836 47874 114888 47880
rect 113732 47796 113784 47802
rect 113732 47738 113784 47744
rect 114560 47796 114612 47802
rect 114560 47738 114612 47744
rect 114572 16574 114600 47738
rect 115952 47734 115980 50102
rect 116032 47864 116084 47870
rect 116032 47806 116084 47812
rect 115940 47728 115992 47734
rect 115940 47670 115992 47676
rect 116044 16574 116072 47806
rect 117332 47598 117360 50102
rect 118160 48074 118188 50102
rect 118148 48068 118200 48074
rect 118148 48010 118200 48016
rect 119264 48006 119292 50102
rect 119252 48000 119304 48006
rect 119252 47942 119304 47948
rect 120368 47802 120396 50102
rect 121564 47870 121592 50102
rect 121552 47864 121604 47870
rect 121552 47806 121604 47812
rect 120356 47796 120408 47802
rect 120356 47738 120408 47744
rect 121460 47796 121512 47802
rect 121460 47738 121512 47744
rect 117320 47592 117372 47598
rect 117320 47534 117372 47540
rect 117320 47116 117372 47122
rect 117320 47058 117372 47064
rect 111996 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 116044 16546 116440 16574
rect 111616 3528 111668 3534
rect 111616 3470 111668 3476
rect 110524 3318 110644 3346
rect 110524 480 110552 3318
rect 111628 480 111656 3470
rect 109286 354 109398 480
rect 109144 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 47058
rect 118792 47048 118844 47054
rect 118792 46990 118844 46996
rect 118804 3534 118832 46990
rect 118884 46980 118936 46986
rect 118884 46922 118936 46928
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 118896 3346 118924 46922
rect 121472 16574 121500 47738
rect 122840 47592 122892 47598
rect 122840 47534 122892 47540
rect 122852 16574 122880 47534
rect 122944 47122 122972 50102
rect 123680 50102 123970 50130
rect 124784 50102 125074 50130
rect 125888 50102 126178 50130
rect 126992 50102 127282 50130
rect 128386 50102 128492 50130
rect 122932 47116 122984 47122
rect 122932 47058 122984 47064
rect 123680 46986 123708 50102
rect 124312 47728 124364 47734
rect 124312 47670 124364 47676
rect 123668 46980 123720 46986
rect 123668 46922 123720 46928
rect 124324 16574 124352 47670
rect 124784 47054 124812 50102
rect 125600 47864 125652 47870
rect 125600 47806 125652 47812
rect 124864 47252 124916 47258
rect 124864 47194 124916 47200
rect 124772 47048 124824 47054
rect 124772 46990 124824 46996
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124324 16546 124720 16574
rect 121092 3800 121144 3806
rect 121092 3742 121144 3748
rect 119896 3528 119948 3534
rect 119896 3470 119948 3476
rect 118804 3318 118924 3346
rect 118804 480 118832 3318
rect 119908 480 119936 3470
rect 121104 480 121132 3742
rect 122300 480 122328 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 124876 3806 124904 47194
rect 124864 3800 124916 3806
rect 124864 3742 124916 3748
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 47806
rect 125888 47258 125916 50102
rect 126992 47802 127020 50102
rect 127072 47932 127124 47938
rect 127072 47874 127124 47880
rect 126980 47796 127032 47802
rect 126980 47738 127032 47744
rect 125876 47252 125928 47258
rect 125876 47194 125928 47200
rect 127084 26234 127112 47874
rect 128464 47598 128492 50102
rect 129200 50102 129490 50130
rect 130304 50102 130594 50130
rect 131408 50102 131698 50130
rect 132604 50102 132710 50130
rect 133432 50102 133814 50130
rect 133984 50102 134918 50130
rect 135640 50102 136022 50130
rect 136744 50102 137126 50130
rect 138032 50102 138230 50130
rect 138952 50102 139334 50130
rect 140056 50102 140438 50130
rect 141160 50102 141542 50130
rect 142264 50102 142646 50130
rect 143552 50102 143658 50130
rect 144472 50102 144762 50130
rect 145576 50102 145866 50130
rect 146680 50102 146970 50130
rect 147876 50102 148074 50130
rect 149072 50102 149178 50130
rect 149992 50102 150282 50130
rect 151096 50102 151386 50130
rect 152200 50102 152490 50130
rect 153304 50102 153594 50130
rect 154592 50102 154698 50130
rect 155328 50102 155710 50130
rect 156432 50102 156814 50130
rect 157536 50102 157918 50130
rect 158732 50102 159022 50130
rect 160126 50102 160232 50130
rect 129200 47734 129228 50102
rect 130304 47870 130332 50102
rect 131408 47870 131436 50102
rect 132604 47938 132632 50102
rect 132592 47932 132644 47938
rect 132592 47874 132644 47880
rect 130292 47864 130344 47870
rect 130292 47806 130344 47812
rect 130476 47864 130528 47870
rect 130476 47806 130528 47812
rect 131396 47864 131448 47870
rect 131396 47806 131448 47812
rect 129188 47728 129240 47734
rect 129188 47670 129240 47676
rect 128452 47592 128504 47598
rect 128452 47534 128504 47540
rect 130384 47048 130436 47054
rect 130384 46990 130436 46996
rect 126992 26206 127112 26234
rect 126992 3534 127020 26206
rect 130396 3534 130424 46990
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 126980 3392 127032 3398
rect 126980 3334 127032 3340
rect 126992 480 127020 3334
rect 128188 480 128216 3470
rect 129384 480 129412 3470
rect 130488 3398 130516 47806
rect 132592 47728 132644 47734
rect 132592 47670 132644 47676
rect 131212 47660 131264 47666
rect 131212 47602 131264 47608
rect 131224 26234 131252 47602
rect 132604 26234 132632 47670
rect 133432 47054 133460 50102
rect 133880 47864 133932 47870
rect 133880 47806 133932 47812
rect 133420 47048 133472 47054
rect 133420 46990 133472 46996
rect 131132 26206 131252 26234
rect 132512 26206 132632 26234
rect 131132 16574 131160 26206
rect 132512 16574 132540 26206
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 130568 3596 130620 3602
rect 130568 3538 130620 3544
rect 130476 3392 130528 3398
rect 130476 3334 130528 3340
rect 130580 480 130608 3538
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 47806
rect 133984 3602 134012 50102
rect 135640 47666 135668 50102
rect 136640 47796 136692 47802
rect 136640 47738 136692 47744
rect 135628 47660 135680 47666
rect 135628 47602 135680 47608
rect 135444 47388 135496 47394
rect 135444 47330 135496 47336
rect 135456 6914 135484 47330
rect 136652 16574 136680 47738
rect 136744 47734 136772 50102
rect 138032 47870 138060 50102
rect 138020 47864 138072 47870
rect 138020 47806 138072 47812
rect 136732 47728 136784 47734
rect 136732 47670 136784 47676
rect 137284 47660 137336 47666
rect 137284 47602 137336 47608
rect 136652 16546 137232 16574
rect 135272 6886 135484 6914
rect 133972 3596 134024 3602
rect 133972 3538 134024 3544
rect 135272 480 135300 6886
rect 136456 3188 136508 3194
rect 136456 3130 136508 3136
rect 136468 480 136496 3130
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 3194 137324 47602
rect 138952 47394 138980 50102
rect 140056 47666 140084 50102
rect 141160 47802 141188 50102
rect 141148 47796 141200 47802
rect 141148 47738 141200 47744
rect 140044 47660 140096 47666
rect 140044 47602 140096 47608
rect 142160 47524 142212 47530
rect 142160 47466 142212 47472
rect 138940 47388 138992 47394
rect 138940 47330 138992 47336
rect 139492 47048 139544 47054
rect 139492 46990 139544 46996
rect 139504 26234 139532 46990
rect 140872 46980 140924 46986
rect 140872 46922 140924 46928
rect 139412 26206 139532 26234
rect 139412 16574 139440 26206
rect 140884 16574 140912 46922
rect 139412 16546 139624 16574
rect 140884 16546 141280 16574
rect 138848 3596 138900 3602
rect 138848 3538 138900 3544
rect 137284 3188 137336 3194
rect 137284 3130 137336 3136
rect 138860 480 138888 3538
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 47466
rect 142264 3602 142292 50102
rect 143552 47054 143580 50102
rect 143816 47864 143868 47870
rect 143816 47806 143868 47812
rect 143632 47592 143684 47598
rect 143632 47534 143684 47540
rect 143540 47048 143592 47054
rect 143540 46990 143592 46996
rect 143644 3602 143672 47534
rect 143828 6914 143856 47806
rect 144472 46986 144500 50102
rect 144920 47932 144972 47938
rect 144920 47874 144972 47880
rect 144460 46980 144512 46986
rect 144460 46922 144512 46928
rect 144932 16574 144960 47874
rect 145576 47530 145604 50102
rect 146680 47870 146708 50102
rect 146668 47864 146720 47870
rect 146668 47806 146720 47812
rect 146300 47796 146352 47802
rect 146300 47738 146352 47744
rect 145564 47524 145616 47530
rect 145564 47466 145616 47472
rect 146312 16574 146340 47738
rect 147772 47660 147824 47666
rect 147772 47602 147824 47608
rect 147784 16574 147812 47602
rect 147876 47598 147904 50102
rect 149072 47938 149100 50102
rect 149060 47932 149112 47938
rect 149060 47874 149112 47880
rect 149992 47802 150020 50102
rect 149980 47796 150032 47802
rect 149980 47738 150032 47744
rect 151096 47666 151124 50102
rect 151820 47932 151872 47938
rect 151820 47874 151872 47880
rect 151084 47660 151136 47666
rect 151084 47602 151136 47608
rect 147864 47592 147916 47598
rect 147864 47534 147916 47540
rect 150532 47048 150584 47054
rect 150532 46990 150584 46996
rect 149244 46980 149296 46986
rect 149244 46922 149296 46928
rect 149256 16574 149284 46922
rect 150544 26234 150572 46990
rect 150452 26206 150572 26234
rect 150452 16574 150480 26206
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147784 16546 147904 16574
rect 149256 16546 149560 16574
rect 150452 16546 150664 16574
rect 143736 6886 143856 6914
rect 142252 3596 142304 3602
rect 142252 3538 142304 3544
rect 143632 3596 143684 3602
rect 143632 3538 143684 3544
rect 143736 3482 143764 6886
rect 144736 3596 144788 3602
rect 144736 3538 144788 3544
rect 143552 3454 143764 3482
rect 143552 480 143580 3454
rect 144748 480 144776 3538
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 9674 151860 47874
rect 151912 47728 151964 47734
rect 151912 47670 151964 47676
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 47670
rect 152200 46986 152228 50102
rect 153304 47054 153332 50102
rect 153384 47864 153436 47870
rect 153384 47806 153436 47812
rect 153292 47048 153344 47054
rect 153292 46990 153344 46996
rect 152188 46980 152240 46986
rect 152188 46922 152240 46928
rect 153396 45554 153424 47806
rect 154592 47734 154620 50102
rect 155328 47938 155356 50102
rect 155316 47932 155368 47938
rect 155316 47874 155368 47880
rect 156432 47870 156460 50102
rect 156420 47864 156472 47870
rect 156420 47806 156472 47812
rect 157432 47864 157484 47870
rect 157432 47806 157484 47812
rect 154580 47728 154632 47734
rect 154580 47670 154632 47676
rect 154580 47592 154632 47598
rect 154580 47534 154632 47540
rect 153304 45526 153424 45554
rect 153304 16574 153332 45526
rect 154592 16574 154620 47534
rect 156052 47524 156104 47530
rect 156052 47466 156104 47472
rect 156064 16574 156092 47466
rect 157444 16574 157472 47806
rect 157536 47598 157564 50102
rect 157524 47592 157576 47598
rect 157524 47534 157576 47540
rect 158732 47530 158760 50102
rect 160204 47870 160232 50102
rect 160848 50102 161230 50130
rect 161952 50102 162334 50130
rect 163056 50102 163438 50130
rect 164252 50102 164542 50130
rect 165540 50102 165646 50130
rect 165724 50102 166750 50130
rect 167472 50102 167762 50130
rect 168484 50102 168866 50130
rect 169772 50102 169970 50130
rect 170048 50102 171074 50130
rect 171888 50102 172178 50130
rect 172624 50102 173282 50130
rect 174096 50102 174386 50130
rect 175292 50102 175490 50130
rect 175568 50102 176594 50130
rect 176672 50102 177698 50130
rect 178052 50102 178802 50130
rect 179524 50102 179814 50130
rect 180812 50102 180918 50130
rect 180996 50102 182022 50130
rect 182192 50102 183126 50130
rect 183572 50102 184230 50130
rect 184952 50102 185334 50130
rect 186438 50102 186544 50130
rect 160192 47864 160244 47870
rect 160192 47806 160244 47812
rect 160848 47666 160876 50102
rect 161572 47932 161624 47938
rect 161572 47874 161624 47880
rect 158812 47660 158864 47666
rect 158812 47602 158864 47608
rect 160836 47660 160888 47666
rect 160836 47602 160888 47608
rect 158720 47524 158772 47530
rect 158720 47466 158772 47472
rect 158824 16574 158852 47602
rect 160100 47048 160152 47054
rect 160100 46990 160152 46996
rect 153304 16546 153792 16574
rect 154592 16546 155448 16574
rect 156064 16546 156184 16574
rect 157444 16546 157840 16574
rect 158824 16546 158944 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 11762 160140 46990
rect 160284 46980 160336 46986
rect 160284 46922 160336 46928
rect 160296 26234 160324 46922
rect 161584 26234 161612 47874
rect 161952 46986 161980 50102
rect 162952 47660 163004 47666
rect 162952 47602 163004 47608
rect 161940 46980 161992 46986
rect 161940 46922 161992 46928
rect 160204 26206 160324 26234
rect 161492 26206 161612 26234
rect 160100 11756 160152 11762
rect 160100 11698 160152 11704
rect 160204 6914 160232 26206
rect 161492 16574 161520 26206
rect 162964 16574 162992 47602
rect 163056 47054 163084 50102
rect 164252 47938 164280 50102
rect 165540 49858 165568 50102
rect 165540 49830 165660 49858
rect 164240 47932 164292 47938
rect 164240 47874 164292 47880
rect 165632 47666 165660 49830
rect 165620 47660 165672 47666
rect 165620 47602 165672 47608
rect 165620 47388 165672 47394
rect 165620 47330 165672 47336
rect 163044 47048 163096 47054
rect 163044 46990 163096 46996
rect 161492 16546 162072 16574
rect 162964 16546 163728 16574
rect 161296 11756 161348 11762
rect 161296 11698 161348 11704
rect 160112 6886 160232 6914
rect 160112 480 160140 6886
rect 161308 480 161336 11698
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 164884 3052 164936 3058
rect 164884 2994 164936 3000
rect 164896 480 164924 2994
rect 165632 1306 165660 47330
rect 165724 3058 165752 50102
rect 167472 47394 167500 50102
rect 168380 47660 168432 47666
rect 168380 47602 168432 47608
rect 167460 47388 167512 47394
rect 167460 47330 167512 47336
rect 165712 3052 165764 3058
rect 165712 2994 165764 3000
rect 167184 3052 167236 3058
rect 167184 2994 167236 3000
rect 165632 1278 166120 1306
rect 166092 480 166120 1278
rect 167196 480 167224 2994
rect 168392 480 168420 47602
rect 168484 3058 168512 50102
rect 169772 47666 169800 50102
rect 169760 47660 169812 47666
rect 169760 47602 169812 47608
rect 169760 46980 169812 46986
rect 169760 46922 169812 46928
rect 169772 3534 169800 46922
rect 170048 45554 170076 50102
rect 171888 46986 171916 50102
rect 172520 47252 172572 47258
rect 172520 47194 172572 47200
rect 171876 46980 171928 46986
rect 171876 46922 171928 46928
rect 169864 45526 170076 45554
rect 169760 3528 169812 3534
rect 169760 3470 169812 3476
rect 169864 3346 169892 45526
rect 172532 3534 172560 47194
rect 170404 3528 170456 3534
rect 170404 3470 170456 3476
rect 172520 3528 172572 3534
rect 172520 3470 172572 3476
rect 169588 3318 169892 3346
rect 168472 3052 168524 3058
rect 168472 2994 168524 3000
rect 169588 480 169616 3318
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170416 354 170444 3470
rect 172624 2802 172652 50102
rect 173900 47796 173952 47802
rect 173900 47738 173952 47744
rect 172796 3528 172848 3534
rect 172796 3470 172848 3476
rect 172440 2774 172652 2802
rect 170742 354 170854 480
rect 170416 326 170854 354
rect 170742 -960 170854 326
rect 171938 354 172050 480
rect 172440 354 172468 2774
rect 171938 326 172468 354
rect 172808 354 172836 3470
rect 173134 354 173246 480
rect 172808 326 173246 354
rect 173912 354 173940 47738
rect 174096 47258 174124 50102
rect 175292 47802 175320 50102
rect 175280 47796 175332 47802
rect 175280 47738 175332 47744
rect 174084 47252 174136 47258
rect 174084 47194 174136 47200
rect 175568 45554 175596 50102
rect 175384 45526 175596 45554
rect 175384 16574 175412 45526
rect 175384 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 480 176700 50102
rect 178052 3482 178080 50102
rect 179420 46980 179472 46986
rect 179420 46922 179472 46928
rect 177868 3454 178080 3482
rect 179052 3528 179104 3534
rect 179052 3470 179104 3476
rect 177868 480 177896 3454
rect 179064 480 179092 3470
rect 179432 3346 179460 46922
rect 179524 3534 179552 50102
rect 180812 46986 180840 50102
rect 180800 46980 180852 46986
rect 180800 46922 180852 46928
rect 179512 3528 179564 3534
rect 179512 3470 179564 3476
rect 179432 3318 180288 3346
rect 180260 480 180288 3318
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 171938 -960 172050 326
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 50102
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 50102
rect 183572 16574 183600 50102
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 480 184980 50102
rect 186320 47864 186372 47870
rect 186320 47806 186372 47812
rect 186332 3534 186360 47806
rect 186516 45554 186544 50102
rect 187160 50102 187542 50130
rect 187712 50102 188646 50130
rect 189092 50102 189750 50130
rect 190472 50102 190762 50130
rect 191866 50102 191972 50130
rect 187160 47870 187188 50102
rect 187148 47864 187200 47870
rect 187148 47806 187200 47812
rect 186424 45526 186544 45554
rect 186320 3528 186372 3534
rect 186320 3470 186372 3476
rect 186424 3346 186452 45526
rect 187712 16574 187740 50102
rect 189092 16574 189120 50102
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186964 3528 187016 3534
rect 186964 3470 187016 3476
rect 186148 3318 186452 3346
rect 186148 480 186176 3318
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186976 354 187004 3470
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186976 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 50102
rect 191944 47818 191972 50102
rect 191852 47790 191972 47818
rect 192036 50102 192970 50130
rect 193324 50102 194074 50130
rect 194612 50102 195178 50130
rect 195992 50102 196282 50130
rect 197386 50102 197492 50130
rect 191852 3482 191880 47790
rect 192036 45554 192064 50102
rect 191944 45526 192064 45554
rect 191944 3602 191972 45526
rect 193324 16574 193352 50102
rect 194612 16574 194640 50102
rect 195992 16574 196020 50102
rect 197464 47818 197492 50102
rect 197372 47790 197492 47818
rect 197556 50102 198490 50130
rect 199594 50102 199976 50130
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 191932 3596 191984 3602
rect 191932 3538 191984 3544
rect 193220 3596 193272 3602
rect 193220 3538 193272 3544
rect 191852 3454 192064 3482
rect 192036 480 192064 3454
rect 193232 480 193260 3538
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197372 3482 197400 47790
rect 197556 45554 197584 50102
rect 199948 48142 199976 50102
rect 200224 50102 200698 50130
rect 201696 50102 201802 50130
rect 202432 50102 202814 50130
rect 203918 50102 204208 50130
rect 199936 48136 199988 48142
rect 199936 48078 199988 48084
rect 200120 48136 200172 48142
rect 200120 48078 200172 48084
rect 197464 45526 197584 45554
rect 197464 3602 197492 45526
rect 197452 3596 197504 3602
rect 197452 3538 197504 3544
rect 199108 3596 199160 3602
rect 199108 3538 199160 3544
rect 197372 3454 197952 3482
rect 197924 480 197952 3454
rect 199120 480 199148 3538
rect 200132 3482 200160 48078
rect 200224 3602 200252 50102
rect 201592 47864 201644 47870
rect 201592 47806 201644 47812
rect 200212 3596 200264 3602
rect 200212 3538 200264 3544
rect 201500 3596 201552 3602
rect 201500 3538 201552 3544
rect 200132 3454 200344 3482
rect 200316 480 200344 3454
rect 201512 480 201540 3538
rect 201604 3194 201632 47806
rect 201696 16574 201724 50102
rect 202432 47870 202460 50102
rect 202420 47864 202472 47870
rect 202420 47806 202472 47812
rect 204180 47818 204208 50102
rect 204364 50102 205022 50130
rect 205652 50102 206126 50130
rect 207230 50102 207520 50130
rect 204180 47790 204300 47818
rect 201696 16546 202736 16574
rect 201592 3188 201644 3194
rect 201592 3130 201644 3136
rect 202708 480 202736 16546
rect 204272 3482 204300 47790
rect 204364 3602 204392 50102
rect 204352 3596 204404 3602
rect 204352 3538 204404 3544
rect 205652 3534 205680 50102
rect 207492 47462 207520 50102
rect 207676 50102 208334 50130
rect 208504 50102 209438 50130
rect 209792 50102 210542 50130
rect 211646 50102 211936 50130
rect 212750 50102 213040 50130
rect 207480 47456 207532 47462
rect 207480 47398 207532 47404
rect 207676 45554 207704 50102
rect 208400 47456 208452 47462
rect 208400 47398 208452 47404
rect 207032 45526 207704 45554
rect 207032 3602 207060 45526
rect 206192 3596 206244 3602
rect 206192 3538 206244 3544
rect 207020 3596 207072 3602
rect 207020 3538 207072 3544
rect 205640 3528 205692 3534
rect 204272 3454 205128 3482
rect 205640 3470 205692 3476
rect 203892 3188 203944 3194
rect 203892 3130 203944 3136
rect 203904 480 203932 3130
rect 205100 480 205128 3454
rect 206204 480 206232 3538
rect 207388 3528 207440 3534
rect 207388 3470 207440 3476
rect 208412 3482 208440 47398
rect 208504 16574 208532 50102
rect 208504 16546 208716 16574
rect 207400 480 207428 3470
rect 208412 3454 208624 3482
rect 208596 480 208624 3454
rect 208688 3194 208716 16546
rect 209792 3670 209820 50102
rect 211908 47870 211936 50102
rect 213012 47870 213040 50102
rect 213104 50102 213854 50130
rect 214024 50102 214866 50130
rect 215312 50102 215970 50130
rect 216692 50102 217074 50130
rect 218072 50102 218178 50130
rect 219282 50102 219388 50130
rect 211896 47864 211948 47870
rect 211896 47806 211948 47812
rect 212540 47864 212592 47870
rect 212540 47806 212592 47812
rect 213000 47864 213052 47870
rect 213000 47806 213052 47812
rect 209780 3664 209832 3670
rect 209780 3606 209832 3612
rect 212172 3664 212224 3670
rect 212172 3606 212224 3612
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 208676 3188 208728 3194
rect 208676 3130 208728 3136
rect 209792 480 209820 3470
rect 210976 3188 211028 3194
rect 210976 3130 211028 3136
rect 210988 480 211016 3130
rect 212184 480 212212 3606
rect 212552 3482 212580 47806
rect 213104 45554 213132 50102
rect 213920 47864 213972 47870
rect 213920 47806 213972 47812
rect 212644 45526 213132 45554
rect 212644 3670 212672 45526
rect 212632 3664 212684 3670
rect 212632 3606 212684 3612
rect 213932 3482 213960 47806
rect 214024 3602 214052 50102
rect 214012 3596 214064 3602
rect 214012 3538 214064 3544
rect 212552 3454 213408 3482
rect 213932 3454 214512 3482
rect 213380 480 213408 3454
rect 214484 480 214512 3454
rect 215312 3194 215340 50102
rect 215668 3664 215720 3670
rect 215668 3606 215720 3612
rect 215300 3188 215352 3194
rect 215300 3130 215352 3136
rect 215680 480 215708 3606
rect 216692 3534 216720 50102
rect 218072 3602 218100 50102
rect 219360 46986 219388 50102
rect 219452 50102 220386 50130
rect 220832 50102 221490 50130
rect 222212 50102 222594 50130
rect 223698 50102 223804 50130
rect 219348 46980 219400 46986
rect 219348 46922 219400 46928
rect 216864 3596 216916 3602
rect 216864 3538 216916 3544
rect 218060 3596 218112 3602
rect 218060 3538 218112 3544
rect 216680 3528 216732 3534
rect 216680 3470 216732 3476
rect 216876 480 216904 3538
rect 219256 3528 219308 3534
rect 219256 3470 219308 3476
rect 218060 3188 218112 3194
rect 218060 3130 218112 3136
rect 218072 480 218100 3130
rect 219268 480 219296 3470
rect 219452 3398 219480 50102
rect 220084 46980 220136 46986
rect 220084 46922 220136 46928
rect 220096 3534 220124 46922
rect 220452 3596 220504 3602
rect 220452 3538 220504 3544
rect 220084 3528 220136 3534
rect 220084 3470 220136 3476
rect 219440 3392 219492 3398
rect 219440 3334 219492 3340
rect 220464 480 220492 3538
rect 220832 3466 220860 50102
rect 222212 3534 222240 50102
rect 223580 46504 223632 46510
rect 223580 46446 223632 46452
rect 223592 3602 223620 46446
rect 223776 45554 223804 50102
rect 224512 50102 224802 50130
rect 225814 50102 226104 50130
rect 224512 46510 224540 50102
rect 226076 47870 226104 50102
rect 226352 50102 226918 50130
rect 227824 50102 228022 50130
rect 229126 50102 229416 50130
rect 230230 50102 230428 50130
rect 226064 47864 226116 47870
rect 226064 47806 226116 47812
rect 224500 46504 224552 46510
rect 224500 46446 224552 46452
rect 223684 45526 223804 45554
rect 223580 3596 223632 3602
rect 223580 3538 223632 3544
rect 221556 3528 221608 3534
rect 221556 3470 221608 3476
rect 222200 3528 222252 3534
rect 222200 3470 222252 3476
rect 220820 3460 220872 3466
rect 220820 3402 220872 3408
rect 221568 480 221596 3470
rect 222752 3392 222804 3398
rect 222752 3334 222804 3340
rect 222764 480 222792 3334
rect 223684 3330 223712 45526
rect 226352 16574 226380 50102
rect 227720 47864 227772 47870
rect 227720 47806 227772 47812
rect 226352 16546 226472 16574
rect 226444 4078 226472 16546
rect 226432 4072 226484 4078
rect 226432 4014 226484 4020
rect 227536 3596 227588 3602
rect 227536 3538 227588 3544
rect 225144 3528 225196 3534
rect 225144 3470 225196 3476
rect 223948 3460 224000 3466
rect 223948 3402 224000 3408
rect 223672 3324 223724 3330
rect 223672 3266 223724 3272
rect 223960 480 223988 3402
rect 225156 480 225184 3470
rect 226340 3324 226392 3330
rect 226340 3266 226392 3272
rect 226352 480 226380 3266
rect 227548 480 227576 3538
rect 227732 490 227760 47806
rect 227824 3874 227852 50102
rect 229388 47870 229416 50102
rect 230400 47938 230428 50102
rect 230492 50102 231334 50130
rect 231964 50102 232438 50130
rect 233344 50102 233542 50130
rect 234540 50102 234646 50130
rect 234724 50102 235750 50130
rect 236854 50102 237144 50130
rect 230388 47932 230440 47938
rect 230388 47874 230440 47880
rect 229376 47864 229428 47870
rect 229376 47806 229428 47812
rect 229836 4072 229888 4078
rect 229836 4014 229888 4020
rect 227812 3868 227864 3874
rect 227812 3810 227864 3816
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 227732 462 228312 490
rect 229848 480 229876 4014
rect 230492 3058 230520 50102
rect 231860 47864 231912 47870
rect 231860 47806 231912 47812
rect 231032 3868 231084 3874
rect 231032 3810 231084 3816
rect 230480 3052 230532 3058
rect 230480 2994 230532 3000
rect 231044 480 231072 3810
rect 228284 354 228312 462
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 231872 354 231900 47806
rect 231964 3534 231992 50102
rect 233240 47932 233292 47938
rect 233240 47874 233292 47880
rect 231952 3528 232004 3534
rect 231952 3470 232004 3476
rect 233252 3482 233280 47874
rect 233344 3602 233372 50102
rect 234540 49858 234568 50102
rect 234540 49830 234660 49858
rect 234632 47666 234660 49830
rect 234620 47660 234672 47666
rect 234620 47602 234672 47608
rect 234724 4078 234752 50102
rect 237116 47326 237144 50102
rect 237484 50102 237866 50130
rect 238772 50102 238970 50130
rect 239968 50102 240074 50130
rect 240244 50102 241178 50130
rect 241532 50102 242282 50130
rect 243386 50102 243768 50130
rect 237380 47660 237432 47666
rect 237380 47602 237432 47608
rect 237104 47320 237156 47326
rect 237104 47262 237156 47268
rect 234712 4072 234764 4078
rect 234712 4014 234764 4020
rect 233332 3596 233384 3602
rect 233332 3538 233384 3544
rect 237012 3596 237064 3602
rect 237012 3538 237064 3544
rect 235816 3528 235868 3534
rect 233252 3454 233464 3482
rect 235816 3470 235868 3476
rect 233436 480 233464 3454
rect 234620 3052 234672 3058
rect 234620 2994 234672 3000
rect 234632 480 234660 2994
rect 235828 480 235856 3470
rect 237024 480 237052 3538
rect 237392 490 237420 47602
rect 237484 3738 237512 50102
rect 237472 3732 237524 3738
rect 237472 3674 237524 3680
rect 238772 3330 238800 50102
rect 239968 47666 239996 50102
rect 239956 47660 240008 47666
rect 239956 47602 240008 47608
rect 240140 47320 240192 47326
rect 240140 47262 240192 47268
rect 239312 4072 239364 4078
rect 239312 4014 239364 4020
rect 238760 3324 238812 3330
rect 238760 3266 238812 3272
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 237392 462 237696 490
rect 239324 480 239352 4014
rect 237668 354 237696 462
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 47262
rect 240244 3466 240272 50102
rect 240784 47660 240836 47666
rect 240784 47602 240836 47608
rect 240796 3534 240824 47602
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 240232 3460 240284 3466
rect 240232 3402 240284 3408
rect 241532 3398 241560 50102
rect 243740 47666 243768 50102
rect 244384 50102 244490 50130
rect 245304 50102 245594 50130
rect 245672 50102 246698 50130
rect 247052 50102 247802 50130
rect 248432 50102 248906 50130
rect 249812 50102 249918 50130
rect 249996 50102 251022 50130
rect 251192 50102 252126 50130
rect 252572 50102 253230 50130
rect 253952 50102 254334 50130
rect 255438 50102 255544 50130
rect 244280 47864 244332 47870
rect 244280 47806 244332 47812
rect 243728 47660 243780 47666
rect 243728 47602 243780 47608
rect 241704 3732 241756 3738
rect 241704 3674 241756 3680
rect 241520 3392 241572 3398
rect 241520 3334 241572 3340
rect 241716 480 241744 3674
rect 244292 3602 244320 47806
rect 244280 3596 244332 3602
rect 244280 3538 244332 3544
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242900 3324 242952 3330
rect 242900 3266 242952 3272
rect 242912 480 242940 3266
rect 244108 480 244136 3470
rect 244384 2990 244412 50102
rect 245304 47870 245332 50102
rect 245292 47864 245344 47870
rect 245292 47806 245344 47812
rect 245672 3466 245700 50102
rect 246304 47660 246356 47666
rect 246304 47602 246356 47608
rect 246316 3534 246344 47602
rect 247052 3874 247080 50102
rect 247040 3868 247092 3874
rect 247040 3810 247092 3816
rect 246304 3528 246356 3534
rect 246304 3470 246356 3476
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 245200 3460 245252 3466
rect 245200 3402 245252 3408
rect 245660 3460 245712 3466
rect 245660 3402 245712 3408
rect 244372 2984 244424 2990
rect 244372 2926 244424 2932
rect 245212 480 245240 3402
rect 246396 3392 246448 3398
rect 246396 3334 246448 3340
rect 246408 480 246436 3334
rect 247604 480 247632 3470
rect 248432 3398 248460 50102
rect 249812 3534 249840 50102
rect 249996 3738 250024 50102
rect 249984 3732 250036 3738
rect 249984 3674 250036 3680
rect 251192 3602 251220 50102
rect 252572 4146 252600 50102
rect 252560 4140 252612 4146
rect 252560 4082 252612 4088
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 249984 3596 250036 3602
rect 249984 3538 250036 3544
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 249800 3528 249852 3534
rect 249800 3470 249852 3476
rect 248420 3392 248472 3398
rect 248420 3334 248472 3340
rect 248788 2984 248840 2990
rect 248788 2926 248840 2932
rect 248800 480 248828 2926
rect 249996 480 250024 3538
rect 251180 3460 251232 3466
rect 251180 3402 251232 3408
rect 251192 480 251220 3402
rect 252388 480 252416 3810
rect 253480 3392 253532 3398
rect 253480 3334 253532 3340
rect 253492 480 253520 3334
rect 253952 3330 253980 50102
rect 255320 47864 255372 47870
rect 255320 47806 255372 47812
rect 255332 3534 255360 47806
rect 255516 45554 255544 50102
rect 256160 50102 256542 50130
rect 256712 50102 257646 50130
rect 258092 50102 258750 50130
rect 259472 50102 259854 50130
rect 260852 50102 260958 50130
rect 261970 50102 262168 50130
rect 256160 47870 256188 50102
rect 256148 47864 256200 47870
rect 256148 47806 256200 47812
rect 255424 45526 255544 45554
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 255320 3528 255372 3534
rect 255320 3470 255372 3476
rect 253940 3324 253992 3330
rect 253940 3266 253992 3272
rect 254688 480 254716 3470
rect 255424 3126 255452 45526
rect 256712 3806 256740 50102
rect 256700 3800 256752 3806
rect 256700 3742 256752 3748
rect 255872 3732 255924 3738
rect 255872 3674 255924 3680
rect 255412 3120 255464 3126
rect 255412 3062 255464 3068
rect 255884 480 255912 3674
rect 257068 3596 257120 3602
rect 257068 3538 257120 3544
rect 257080 480 257108 3538
rect 258092 3398 258120 50102
rect 258264 4140 258316 4146
rect 258264 4082 258316 4088
rect 258080 3392 258132 3398
rect 258080 3334 258132 3340
rect 258276 480 258304 4082
rect 259472 3602 259500 50102
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 260852 3466 260880 50102
rect 262140 47870 262168 50102
rect 262232 50102 263074 50130
rect 263612 50102 264178 50130
rect 265282 50102 265664 50130
rect 266386 50102 266492 50130
rect 262128 47864 262180 47870
rect 262128 47806 262180 47812
rect 261760 3528 261812 3534
rect 261760 3470 261812 3476
rect 260840 3460 260892 3466
rect 260840 3402 260892 3408
rect 259460 3324 259512 3330
rect 259460 3266 259512 3272
rect 259472 480 259500 3266
rect 260656 3120 260708 3126
rect 260656 3062 260708 3068
rect 260668 480 260696 3062
rect 261772 480 261800 3470
rect 262232 3126 262260 50102
rect 263612 4010 263640 50102
rect 264244 47864 264296 47870
rect 264244 47806 264296 47812
rect 263600 4004 263652 4010
rect 263600 3946 263652 3952
rect 264256 3942 264284 47806
rect 265636 47598 265664 50102
rect 266464 47682 266492 50102
rect 266372 47654 266492 47682
rect 266556 50102 267490 50130
rect 267752 50102 268594 50130
rect 269132 50102 269698 50130
rect 270604 50102 270802 50130
rect 271800 50102 271906 50130
rect 271984 50102 272918 50130
rect 273272 50102 274022 50130
rect 274652 50102 275126 50130
rect 276032 50102 276230 50130
rect 276308 50102 277334 50130
rect 277504 50102 278438 50130
rect 278792 50102 279542 50130
rect 280172 50102 280646 50130
rect 281552 50102 281750 50130
rect 281920 50102 282854 50130
rect 282932 50102 283958 50130
rect 284312 50102 284970 50130
rect 285692 50102 286074 50130
rect 287178 50102 287284 50130
rect 265624 47592 265676 47598
rect 265624 47534 265676 47540
rect 264244 3936 264296 3942
rect 264244 3878 264296 3884
rect 262956 3800 263008 3806
rect 262956 3742 263008 3748
rect 262220 3120 262272 3126
rect 262220 3062 262272 3068
rect 262968 480 262996 3742
rect 266372 3738 266400 47654
rect 266556 45554 266584 50102
rect 266464 45526 266584 45554
rect 266360 3732 266412 3738
rect 266360 3674 266412 3680
rect 266464 3602 266492 45526
rect 267752 16574 267780 50102
rect 267752 16546 267872 16574
rect 267740 3936 267792 3942
rect 267740 3878 267792 3884
rect 265348 3596 265400 3602
rect 265348 3538 265400 3544
rect 266452 3596 266504 3602
rect 266452 3538 266504 3544
rect 264152 3392 264204 3398
rect 264152 3334 264204 3340
rect 264164 480 264192 3334
rect 265360 480 265388 3538
rect 266544 3460 266596 3466
rect 266544 3402 266596 3408
rect 266556 480 266584 3402
rect 267752 480 267780 3878
rect 267844 3398 267872 16546
rect 269132 3466 269160 50102
rect 270500 47592 270552 47598
rect 270500 47534 270552 47540
rect 270040 4004 270092 4010
rect 270040 3946 270092 3952
rect 269120 3460 269172 3466
rect 269120 3402 269172 3408
rect 267832 3392 267884 3398
rect 267832 3334 267884 3340
rect 268844 3120 268896 3126
rect 268844 3062 268896 3068
rect 268856 480 268884 3062
rect 270052 480 270080 3946
rect 270512 490 270540 47534
rect 270604 3534 270632 50102
rect 271800 49858 271828 50102
rect 271800 49830 271920 49858
rect 271892 47870 271920 49830
rect 271880 47864 271932 47870
rect 271880 47806 271932 47812
rect 271984 4078 272012 50102
rect 271972 4072 272024 4078
rect 271972 4014 272024 4020
rect 273272 3738 273300 50102
rect 272432 3732 272484 3738
rect 272432 3674 272484 3680
rect 273260 3732 273312 3738
rect 273260 3674 273312 3680
rect 270592 3528 270644 3534
rect 270592 3470 270644 3476
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270512 462 270816 490
rect 272444 480 272472 3674
rect 274652 3602 274680 50102
rect 276032 3670 276060 50102
rect 276308 45554 276336 50102
rect 277400 47864 277452 47870
rect 277400 47806 277452 47812
rect 276124 45526 276336 45554
rect 276020 3664 276072 3670
rect 276020 3606 276072 3612
rect 273628 3596 273680 3602
rect 273628 3538 273680 3544
rect 274640 3596 274692 3602
rect 274640 3538 274692 3544
rect 273640 480 273668 3538
rect 276124 3466 276152 45526
rect 277124 3528 277176 3534
rect 277412 3516 277440 47806
rect 277504 3942 277532 50102
rect 277492 3936 277544 3942
rect 277492 3878 277544 3884
rect 277412 3488 278360 3516
rect 277124 3470 277176 3476
rect 276020 3460 276072 3466
rect 276020 3402 276072 3408
rect 276112 3460 276164 3466
rect 276112 3402 276164 3408
rect 274824 3392 274876 3398
rect 274824 3334 274876 3340
rect 274836 480 274864 3334
rect 276032 480 276060 3402
rect 277136 480 277164 3470
rect 278332 480 278360 3488
rect 278792 3126 278820 50102
rect 279516 4072 279568 4078
rect 279516 4014 279568 4020
rect 278780 3120 278832 3126
rect 278780 3062 278832 3068
rect 279528 480 279556 4014
rect 280172 3194 280200 50102
rect 280712 3732 280764 3738
rect 280712 3674 280764 3680
rect 280160 3188 280212 3194
rect 280160 3130 280212 3136
rect 280724 480 280752 3674
rect 281552 2990 281580 50102
rect 281920 45554 281948 50102
rect 281644 45526 281948 45554
rect 281644 3874 281672 45526
rect 281632 3868 281684 3874
rect 281632 3810 281684 3816
rect 282932 3806 282960 50102
rect 282920 3800 282972 3806
rect 282920 3742 282972 3748
rect 284312 3670 284340 50102
rect 285692 3942 285720 50102
rect 287060 47864 287112 47870
rect 287060 47806 287112 47812
rect 285404 3936 285456 3942
rect 285404 3878 285456 3884
rect 285680 3936 285732 3942
rect 285680 3878 285732 3884
rect 283104 3664 283156 3670
rect 283104 3606 283156 3612
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 281908 3596 281960 3602
rect 281908 3538 281960 3544
rect 281540 2984 281592 2990
rect 281540 2926 281592 2932
rect 281920 480 281948 3538
rect 283116 480 283144 3606
rect 284300 3460 284352 3466
rect 284300 3402 284352 3408
rect 284312 480 284340 3402
rect 285416 480 285444 3878
rect 286600 3120 286652 3126
rect 286600 3062 286652 3068
rect 286612 480 286640 3062
rect 287072 2922 287100 47806
rect 287256 45554 287284 50102
rect 287992 50102 288282 50130
rect 288452 50102 289386 50130
rect 289832 50102 290490 50130
rect 291212 50102 291594 50130
rect 292592 50102 292698 50130
rect 293802 50102 293908 50130
rect 287992 47870 288020 50102
rect 287980 47864 288032 47870
rect 287980 47806 288032 47812
rect 287164 45526 287284 45554
rect 287164 3602 287192 45526
rect 287152 3596 287204 3602
rect 287152 3538 287204 3544
rect 288452 3466 288480 50102
rect 288440 3460 288492 3466
rect 288440 3402 288492 3408
rect 287796 3188 287848 3194
rect 287796 3130 287848 3136
rect 287060 2916 287112 2922
rect 287060 2858 287112 2864
rect 287808 480 287836 3130
rect 289832 3058 289860 50102
rect 290188 3868 290240 3874
rect 290188 3810 290240 3816
rect 289820 3052 289872 3058
rect 289820 2994 289872 3000
rect 288992 2984 289044 2990
rect 288992 2926 289044 2932
rect 289004 480 289032 2926
rect 290200 480 290228 3810
rect 291212 3534 291240 50102
rect 292592 4146 292620 50102
rect 293880 47598 293908 50102
rect 293972 50102 294906 50130
rect 295352 50102 296010 50130
rect 296732 50102 297022 50130
rect 298126 50102 298232 50130
rect 293868 47592 293920 47598
rect 293868 47534 293920 47540
rect 292580 4140 292632 4146
rect 292580 4082 292632 4088
rect 293684 3936 293736 3942
rect 293684 3878 293736 3884
rect 291384 3800 291436 3806
rect 291384 3742 291436 3748
rect 291200 3528 291252 3534
rect 291200 3470 291252 3476
rect 291396 480 291424 3742
rect 292580 3664 292632 3670
rect 292580 3606 292632 3612
rect 292592 480 292620 3606
rect 293696 480 293724 3878
rect 293972 3670 294000 50102
rect 295352 4078 295380 50102
rect 295340 4072 295392 4078
rect 295340 4014 295392 4020
rect 293960 3664 294012 3670
rect 293960 3606 294012 3612
rect 294880 3596 294932 3602
rect 294880 3538 294932 3544
rect 294892 480 294920 3538
rect 296732 3330 296760 50102
rect 298204 47818 298232 50102
rect 298112 47790 298232 47818
rect 298388 50102 299230 50130
rect 299492 50102 300334 50130
rect 300872 50102 301438 50130
rect 302252 50102 302542 50130
rect 303646 50102 303752 50130
rect 298112 4010 298140 47790
rect 298388 45554 298416 50102
rect 298204 45526 298416 45554
rect 298100 4004 298152 4010
rect 298100 3946 298152 3952
rect 298204 3466 298232 45526
rect 299492 3806 299520 50102
rect 300124 47592 300176 47598
rect 300124 47534 300176 47540
rect 299480 3800 299532 3806
rect 299480 3742 299532 3748
rect 299664 3528 299716 3534
rect 299664 3470 299716 3476
rect 297272 3460 297324 3466
rect 297272 3402 297324 3408
rect 298192 3460 298244 3466
rect 298192 3402 298244 3408
rect 296720 3324 296772 3330
rect 296720 3266 296772 3272
rect 296076 2916 296128 2922
rect 296076 2858 296128 2864
rect 296088 480 296116 2858
rect 297284 480 297312 3402
rect 298468 3052 298520 3058
rect 298468 2994 298520 3000
rect 298480 480 298508 2994
rect 299676 480 299704 3470
rect 300136 3058 300164 47534
rect 300768 4140 300820 4146
rect 300768 4082 300820 4088
rect 300124 3052 300176 3058
rect 300124 2994 300176 3000
rect 300780 480 300808 4082
rect 300872 3398 300900 50102
rect 302252 4146 302280 50102
rect 303724 47818 303752 50102
rect 303632 47790 303752 47818
rect 303816 50102 304750 50130
rect 305012 50102 305854 50130
rect 306392 50102 306958 50130
rect 307970 50102 308076 50130
rect 302240 4140 302292 4146
rect 302240 4082 302292 4088
rect 303632 3942 303660 47790
rect 303816 45554 303844 50102
rect 303724 45526 303844 45554
rect 303620 3936 303672 3942
rect 303620 3878 303672 3884
rect 303160 3664 303212 3670
rect 303160 3606 303212 3612
rect 300860 3392 300912 3398
rect 300860 3334 300912 3340
rect 301964 3052 302016 3058
rect 301964 2994 302016 3000
rect 301976 480 302004 2994
rect 303172 480 303200 3606
rect 303724 3602 303752 45526
rect 304356 4072 304408 4078
rect 304356 4014 304408 4020
rect 303712 3596 303764 3602
rect 303712 3538 303764 3544
rect 304368 480 304396 4014
rect 305012 3738 305040 50102
rect 306392 3874 306420 50102
rect 308048 47870 308076 50102
rect 308140 50102 309074 50130
rect 309152 50102 310178 50130
rect 310532 50102 311282 50130
rect 311912 50102 312386 50130
rect 313384 50102 313490 50130
rect 314304 50102 314594 50130
rect 314672 50102 315698 50130
rect 316052 50102 316802 50130
rect 317432 50102 317906 50130
rect 318812 50102 319010 50130
rect 320022 50102 320128 50130
rect 308036 47864 308088 47870
rect 308036 47806 308088 47812
rect 308140 45554 308168 50102
rect 307772 45526 308168 45554
rect 306748 4004 306800 4010
rect 306748 3946 306800 3952
rect 306380 3868 306432 3874
rect 306380 3810 306432 3816
rect 305000 3732 305052 3738
rect 305000 3674 305052 3680
rect 305552 3324 305604 3330
rect 305552 3266 305604 3272
rect 305564 480 305592 3266
rect 306760 480 306788 3946
rect 307772 3670 307800 45526
rect 309048 3800 309100 3806
rect 309048 3742 309100 3748
rect 307760 3664 307812 3670
rect 307760 3606 307812 3612
rect 307944 3460 307996 3466
rect 307944 3402 307996 3408
rect 307956 480 307984 3402
rect 309060 480 309088 3742
rect 309152 3534 309180 50102
rect 309784 47864 309836 47870
rect 309784 47806 309836 47812
rect 309796 4078 309824 47806
rect 309784 4072 309836 4078
rect 309784 4014 309836 4020
rect 310532 4010 310560 50102
rect 311440 4140 311492 4146
rect 311440 4082 311492 4088
rect 310520 4004 310572 4010
rect 310520 3946 310572 3952
rect 309140 3528 309192 3534
rect 309140 3470 309192 3476
rect 310244 3392 310296 3398
rect 310244 3334 310296 3340
rect 310256 480 310284 3334
rect 311452 480 311480 4082
rect 311912 3806 311940 50102
rect 313280 47864 313332 47870
rect 313280 47806 313332 47812
rect 313292 4146 313320 47806
rect 313280 4140 313332 4146
rect 313280 4082 313332 4088
rect 312636 3936 312688 3942
rect 312636 3878 312688 3884
rect 311900 3800 311952 3806
rect 311900 3742 311952 3748
rect 312648 480 312676 3878
rect 313384 3398 313412 50102
rect 314304 47870 314332 50102
rect 314292 47864 314344 47870
rect 314292 47806 314344 47812
rect 314672 3602 314700 50102
rect 316052 3738 316080 50102
rect 317328 4072 317380 4078
rect 317328 4014 317380 4020
rect 316224 3868 316276 3874
rect 316224 3810 316276 3816
rect 315028 3732 315080 3738
rect 315028 3674 315080 3680
rect 316040 3732 316092 3738
rect 316040 3674 316092 3680
rect 313832 3596 313884 3602
rect 313832 3538 313884 3544
rect 314660 3596 314712 3602
rect 314660 3538 314712 3544
rect 313372 3392 313424 3398
rect 313372 3334 313424 3340
rect 313844 480 313872 3538
rect 315040 480 315068 3674
rect 316236 480 316264 3810
rect 317340 480 317368 4014
rect 317432 3874 317460 50102
rect 318812 3942 318840 50102
rect 320100 47870 320128 50102
rect 320192 50102 321126 50130
rect 321572 50102 322230 50130
rect 322952 50102 323334 50130
rect 324332 50102 324438 50130
rect 324516 50102 325542 50130
rect 325712 50102 326646 50130
rect 327092 50102 327750 50130
rect 328472 50102 328854 50130
rect 329958 50102 330064 50130
rect 320088 47864 320140 47870
rect 320088 47806 320140 47812
rect 318800 3936 318852 3942
rect 318800 3878 318852 3884
rect 317420 3868 317472 3874
rect 317420 3810 317472 3816
rect 320192 3670 320220 50102
rect 320916 4004 320968 4010
rect 320916 3946 320968 3952
rect 318524 3664 318576 3670
rect 318524 3606 318576 3612
rect 320180 3664 320232 3670
rect 320180 3606 320232 3612
rect 318536 480 318564 3606
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 319732 480 319760 3470
rect 320928 480 320956 3946
rect 321572 3534 321600 50102
rect 322952 4078 322980 50102
rect 323584 47864 323636 47870
rect 323584 47806 323636 47812
rect 322940 4072 322992 4078
rect 322940 4014 322992 4020
rect 323596 4010 323624 47806
rect 323584 4004 323636 4010
rect 323584 3946 323636 3952
rect 322112 3800 322164 3806
rect 322112 3742 322164 3748
rect 321560 3528 321612 3534
rect 321560 3470 321612 3476
rect 322124 480 322152 3742
rect 323308 3392 323360 3398
rect 323308 3334 323360 3340
rect 323320 480 323348 3334
rect 324332 3194 324360 50102
rect 324412 4140 324464 4146
rect 324412 4082 324464 4088
rect 324320 3188 324372 3194
rect 324320 3130 324372 3136
rect 324424 480 324452 4082
rect 324516 3466 324544 50102
rect 325712 3602 325740 50102
rect 327092 3738 327120 50102
rect 328000 3868 328052 3874
rect 328000 3810 328052 3816
rect 326804 3732 326856 3738
rect 326804 3674 326856 3680
rect 327080 3732 327132 3738
rect 327080 3674 327132 3680
rect 325608 3596 325660 3602
rect 325608 3538 325660 3544
rect 325700 3596 325752 3602
rect 325700 3538 325752 3544
rect 324504 3460 324556 3466
rect 324504 3402 324556 3408
rect 325620 480 325648 3538
rect 326816 480 326844 3674
rect 328012 480 328040 3810
rect 328472 3806 328500 50102
rect 329840 47864 329892 47870
rect 329840 47806 329892 47812
rect 329196 3936 329248 3942
rect 329196 3878 329248 3884
rect 328460 3800 328512 3806
rect 328460 3742 328512 3748
rect 329208 480 329236 3878
rect 329852 3874 329880 47806
rect 330036 45554 330064 50102
rect 330680 50102 331062 50130
rect 331232 50102 332074 50130
rect 332612 50102 333178 50130
rect 333992 50102 334282 50130
rect 335386 50102 335492 50130
rect 330680 47870 330708 50102
rect 330668 47864 330720 47870
rect 330668 47806 330720 47812
rect 329944 45526 330064 45554
rect 329840 3868 329892 3874
rect 329840 3810 329892 3816
rect 329944 3262 329972 45526
rect 330392 4004 330444 4010
rect 330392 3946 330444 3952
rect 329932 3256 329984 3262
rect 329932 3198 329984 3204
rect 330404 480 330432 3946
rect 331232 3330 331260 50102
rect 332612 3942 332640 50102
rect 333992 4078 334020 50102
rect 335464 47818 335492 50102
rect 335372 47790 335492 47818
rect 335556 50102 336490 50130
rect 336752 50102 337594 50130
rect 338132 50102 338698 50130
rect 339512 50102 339802 50130
rect 340906 50102 341012 50130
rect 333888 4072 333940 4078
rect 333888 4014 333940 4020
rect 333980 4072 334032 4078
rect 333980 4014 334032 4020
rect 332600 3936 332652 3942
rect 332600 3878 332652 3884
rect 331588 3664 331640 3670
rect 331588 3606 331640 3612
rect 331220 3324 331272 3330
rect 331220 3266 331272 3272
rect 331600 480 331628 3606
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 332704 480 332732 3470
rect 333900 480 333928 4014
rect 335372 3670 335400 47790
rect 335556 45554 335584 50102
rect 335464 45526 335584 45554
rect 335360 3664 335412 3670
rect 335360 3606 335412 3612
rect 335464 3534 335492 45526
rect 335452 3528 335504 3534
rect 335452 3470 335504 3476
rect 336752 3466 336780 50102
rect 338132 4010 338160 50102
rect 339512 4146 339540 50102
rect 340984 47682 341012 50102
rect 340892 47654 341012 47682
rect 341076 50102 342010 50130
rect 342272 50102 343114 50130
rect 343652 50102 344126 50130
rect 345032 50102 345230 50130
rect 345308 50102 346334 50130
rect 347438 50102 347728 50130
rect 339500 4140 339552 4146
rect 339500 4082 339552 4088
rect 338120 4004 338172 4010
rect 338120 3946 338172 3952
rect 339868 3800 339920 3806
rect 339868 3742 339920 3748
rect 338672 3732 338724 3738
rect 338672 3674 338724 3680
rect 337476 3596 337528 3602
rect 337476 3538 337528 3544
rect 336280 3460 336332 3466
rect 336280 3402 336332 3408
rect 336740 3460 336792 3466
rect 336740 3402 336792 3408
rect 335084 3188 335136 3194
rect 335084 3130 335136 3136
rect 335096 480 335124 3130
rect 336292 480 336320 3402
rect 337488 480 337516 3538
rect 338684 480 338712 3674
rect 339880 480 339908 3742
rect 340892 3398 340920 47654
rect 341076 45554 341104 50102
rect 340984 45526 341104 45554
rect 340984 16574 341012 45526
rect 340984 16546 341104 16574
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 341076 3262 341104 16546
rect 342168 3868 342220 3874
rect 342168 3810 342220 3816
rect 340972 3256 341024 3262
rect 340972 3198 341024 3204
rect 341064 3256 341116 3262
rect 341064 3198 341116 3204
rect 340984 480 341012 3198
rect 342180 480 342208 3810
rect 342272 3602 342300 50102
rect 343652 3806 343680 50102
rect 345032 3942 345060 50102
rect 345308 45554 345336 50102
rect 347700 47598 347728 50102
rect 347792 50102 348542 50130
rect 349172 50102 349646 50130
rect 350644 50102 350750 50130
rect 350828 50102 351854 50130
rect 351932 50102 352958 50130
rect 353312 50102 354062 50130
rect 354692 50102 355074 50130
rect 356072 50102 356178 50130
rect 356256 50102 357282 50130
rect 357452 50102 358386 50130
rect 358832 50102 359490 50130
rect 360212 50102 360594 50130
rect 361698 50102 362080 50130
rect 362802 50102 362908 50130
rect 347688 47592 347740 47598
rect 347688 47534 347740 47540
rect 345124 45526 345336 45554
rect 344560 3936 344612 3942
rect 344560 3878 344612 3884
rect 345020 3936 345072 3942
rect 345020 3878 345072 3884
rect 343640 3800 343692 3806
rect 343640 3742 343692 3748
rect 342260 3596 342312 3602
rect 342260 3538 342312 3544
rect 343364 3324 343416 3330
rect 343364 3266 343416 3272
rect 343376 480 343404 3266
rect 344572 480 344600 3878
rect 345124 3330 345152 45526
rect 347792 4078 347820 50102
rect 345756 4072 345808 4078
rect 345756 4014 345808 4020
rect 347780 4072 347832 4078
rect 347780 4014 347832 4020
rect 345112 3324 345164 3330
rect 345112 3266 345164 3272
rect 345768 480 345796 4014
rect 349172 3738 349200 50102
rect 350644 47666 350672 50102
rect 350632 47660 350684 47666
rect 350632 47602 350684 47608
rect 350828 45554 350856 50102
rect 350552 45526 350856 45554
rect 350448 4004 350500 4010
rect 350448 3946 350500 3952
rect 349160 3732 349212 3738
rect 349160 3674 349212 3680
rect 346952 3664 347004 3670
rect 346952 3606 347004 3612
rect 346964 480 346992 3606
rect 348056 3528 348108 3534
rect 348056 3470 348108 3476
rect 348068 480 348096 3470
rect 349252 3460 349304 3466
rect 349252 3402 349304 3408
rect 349264 480 349292 3402
rect 350460 480 350488 3946
rect 350552 3534 350580 45526
rect 351644 4140 351696 4146
rect 351644 4082 351696 4088
rect 350540 3528 350592 3534
rect 350540 3470 350592 3476
rect 351656 480 351684 4082
rect 351932 3670 351960 50102
rect 351920 3664 351972 3670
rect 351920 3606 351972 3612
rect 353312 3398 353340 50102
rect 354692 3874 354720 50102
rect 356072 4146 356100 50102
rect 356060 4140 356112 4146
rect 356060 4082 356112 4088
rect 356256 4010 356284 50102
rect 356244 4004 356296 4010
rect 356244 3946 356296 3952
rect 354680 3868 354732 3874
rect 354680 3810 354732 3816
rect 357452 3806 357480 50102
rect 358084 47592 358136 47598
rect 358084 47534 358136 47540
rect 357532 3936 357584 3942
rect 357532 3878 357584 3884
rect 356336 3800 356388 3806
rect 356336 3742 356388 3748
rect 357440 3800 357492 3806
rect 357440 3742 357492 3748
rect 355232 3596 355284 3602
rect 355232 3538 355284 3544
rect 352840 3392 352892 3398
rect 352840 3334 352892 3340
rect 353300 3392 353352 3398
rect 353300 3334 353352 3340
rect 352852 480 352880 3334
rect 354036 3256 354088 3262
rect 354036 3198 354088 3204
rect 354048 480 354076 3198
rect 355244 480 355272 3538
rect 356348 480 356376 3742
rect 357544 480 357572 3878
rect 358096 3534 358124 47534
rect 358832 3602 358860 50102
rect 360212 3942 360240 50102
rect 362052 46986 362080 50102
rect 362880 47734 362908 50102
rect 362972 50102 363906 50130
rect 364352 50102 365010 50130
rect 365732 50102 366114 50130
rect 367020 50102 367126 50130
rect 367204 50102 368230 50130
rect 368492 50102 369334 50130
rect 370438 50102 370728 50130
rect 362868 47728 362920 47734
rect 362868 47670 362920 47676
rect 362224 47660 362276 47666
rect 362224 47602 362276 47608
rect 362040 46980 362092 46986
rect 362040 46922 362092 46928
rect 361120 4072 361172 4078
rect 361120 4014 361172 4020
rect 360200 3936 360252 3942
rect 360200 3878 360252 3884
rect 358820 3596 358872 3602
rect 358820 3538 358872 3544
rect 358084 3528 358136 3534
rect 358084 3470 358136 3476
rect 359924 3528 359976 3534
rect 359924 3470 359976 3476
rect 358728 3324 358780 3330
rect 358728 3266 358780 3272
rect 358740 480 358768 3266
rect 359936 480 359964 3470
rect 361132 480 361160 4014
rect 362236 3534 362264 47602
rect 362972 4078 363000 50102
rect 362960 4072 363012 4078
rect 362960 4014 363012 4020
rect 364352 3806 364380 50102
rect 364340 3800 364392 3806
rect 364340 3742 364392 3748
rect 362316 3732 362368 3738
rect 362316 3674 362368 3680
rect 362224 3528 362276 3534
rect 362224 3470 362276 3476
rect 362328 480 362356 3674
rect 365732 3534 365760 50102
rect 367020 49858 367048 50102
rect 367020 49830 367140 49858
rect 367112 47666 367140 49830
rect 367100 47660 367152 47666
rect 367100 47602 367152 47608
rect 366364 46980 366416 46986
rect 366364 46922 366416 46928
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 363512 3528 363564 3534
rect 363512 3470 363564 3476
rect 365720 3528 365772 3534
rect 365720 3470 365772 3476
rect 363524 480 363552 3470
rect 364616 3460 364668 3466
rect 364616 3402 364668 3408
rect 364628 480 364656 3402
rect 365824 480 365852 3606
rect 366376 3466 366404 46922
rect 367204 3738 367232 50102
rect 368492 3874 368520 50102
rect 370700 47870 370728 50102
rect 371252 50102 371542 50130
rect 372646 50102 372936 50130
rect 373750 50102 373856 50130
rect 370688 47864 370740 47870
rect 370688 47806 370740 47812
rect 369400 4140 369452 4146
rect 369400 4082 369452 4088
rect 368204 3868 368256 3874
rect 368204 3810 368256 3816
rect 368480 3868 368532 3874
rect 368480 3810 368532 3816
rect 367192 3732 367244 3738
rect 367192 3674 367244 3680
rect 366364 3460 366416 3466
rect 366364 3402 366416 3408
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 368216 480 368244 3810
rect 369412 480 369440 4082
rect 371252 4010 371280 50102
rect 372908 47938 372936 50102
rect 372896 47932 372948 47938
rect 372896 47874 372948 47880
rect 373828 47598 373856 50102
rect 374012 50102 374854 50130
rect 375484 50102 375958 50130
rect 377062 50102 377352 50130
rect 378166 50102 378272 50130
rect 373816 47592 373868 47598
rect 373816 47534 373868 47540
rect 370596 4004 370648 4010
rect 370596 3946 370648 3952
rect 371240 4004 371292 4010
rect 371240 3946 371292 3952
rect 370608 480 370636 3946
rect 371700 3664 371752 3670
rect 371700 3606 371752 3612
rect 371712 480 371740 3606
rect 374012 3602 374040 50102
rect 375380 47728 375432 47734
rect 375380 47670 375432 47676
rect 374092 3936 374144 3942
rect 374092 3878 374144 3884
rect 372896 3596 372948 3602
rect 372896 3538 372948 3544
rect 374000 3596 374052 3602
rect 374000 3538 374052 3544
rect 372908 480 372936 3538
rect 374104 480 374132 3878
rect 375288 3460 375340 3466
rect 375288 3402 375340 3408
rect 375300 480 375328 3402
rect 375392 626 375420 47670
rect 375484 3670 375512 50102
rect 377324 47802 377352 50102
rect 378244 47852 378272 50102
rect 378152 47824 378272 47852
rect 378520 50102 379178 50130
rect 380282 50102 380664 50130
rect 377312 47796 377364 47802
rect 377312 47738 377364 47744
rect 377680 4072 377732 4078
rect 377680 4014 377732 4020
rect 375472 3664 375524 3670
rect 375472 3606 375524 3612
rect 375392 598 376064 626
rect 270788 354 270816 462
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 598
rect 377692 480 377720 4014
rect 378152 3398 378180 47824
rect 378520 45554 378548 50102
rect 380636 47734 380664 50102
rect 381004 50102 381386 50130
rect 382292 50102 382490 50130
rect 383488 50102 383594 50130
rect 383764 50102 384698 50130
rect 385052 50102 385802 50130
rect 386906 50102 387288 50130
rect 380624 47728 380676 47734
rect 380624 47670 380676 47676
rect 380900 47660 380952 47666
rect 380900 47602 380952 47608
rect 378244 45526 378548 45554
rect 378140 3392 378192 3398
rect 378140 3334 378192 3340
rect 378244 3330 378272 45526
rect 378876 3800 378928 3806
rect 378876 3742 378928 3748
rect 378232 3324 378284 3330
rect 378232 3266 378284 3272
rect 378888 480 378916 3742
rect 379980 3528 380032 3534
rect 379980 3470 380032 3476
rect 380912 3482 380940 47602
rect 381004 4146 381032 50102
rect 380992 4140 381044 4146
rect 380992 4082 381044 4088
rect 379992 480 380020 3470
rect 380912 3454 381216 3482
rect 382292 3466 382320 50102
rect 383488 47666 383516 50102
rect 383660 47864 383712 47870
rect 383660 47806 383712 47812
rect 383476 47660 383528 47666
rect 383476 47602 383528 47608
rect 383568 3868 383620 3874
rect 383568 3810 383620 3816
rect 382372 3732 382424 3738
rect 382372 3674 382424 3680
rect 381188 480 381216 3454
rect 382280 3460 382332 3466
rect 382280 3402 382332 3408
rect 382384 480 382412 3674
rect 383580 480 383608 3810
rect 383672 626 383700 47806
rect 383764 3942 383792 50102
rect 383752 3936 383804 3942
rect 383752 3878 383804 3884
rect 385052 3738 385080 50102
rect 385684 47932 385736 47938
rect 385684 47874 385736 47880
rect 385040 3732 385092 3738
rect 385040 3674 385092 3680
rect 385696 3534 385724 47874
rect 387260 47870 387288 50102
rect 387904 50102 388010 50130
rect 388088 50102 389114 50130
rect 390126 50102 390416 50130
rect 387248 47864 387300 47870
rect 387248 47806 387300 47812
rect 387800 47592 387852 47598
rect 387800 47534 387852 47540
rect 385960 4004 386012 4010
rect 385960 3946 386012 3952
rect 385684 3528 385736 3534
rect 385684 3470 385736 3476
rect 383672 598 384344 626
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 598
rect 385972 480 386000 3946
rect 387156 3528 387208 3534
rect 387156 3470 387208 3476
rect 387168 480 387196 3470
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 47534
rect 387904 4078 387932 50102
rect 387892 4072 387944 4078
rect 387892 4014 387944 4020
rect 388088 3534 388116 50102
rect 390388 47598 390416 50102
rect 390664 50102 391230 50130
rect 391952 50102 392334 50130
rect 393332 50102 393438 50130
rect 393516 50102 394542 50130
rect 394804 50102 395646 50130
rect 396750 50102 397040 50130
rect 390376 47592 390428 47598
rect 390376 47534 390428 47540
rect 390664 3670 390692 50102
rect 390744 47796 390796 47802
rect 390744 47738 390796 47744
rect 390756 16574 390784 47738
rect 390756 16546 391888 16574
rect 390560 3664 390612 3670
rect 390560 3606 390612 3612
rect 390652 3664 390704 3670
rect 390652 3606 390704 3612
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 388076 3528 388128 3534
rect 388076 3470 388128 3476
rect 389468 480 389496 3538
rect 390572 1850 390600 3606
rect 390572 1822 390692 1850
rect 390664 480 390692 1822
rect 391860 480 391888 16546
rect 391952 4078 391980 50102
rect 393332 47938 393360 50102
rect 393320 47932 393372 47938
rect 393320 47874 393372 47880
rect 393516 45554 393544 50102
rect 394700 47728 394752 47734
rect 394700 47670 394752 47676
rect 393332 45526 393544 45554
rect 391940 4072 391992 4078
rect 391940 4014 391992 4020
rect 393332 3398 393360 45526
rect 393044 3392 393096 3398
rect 393044 3334 393096 3340
rect 393320 3392 393372 3398
rect 393320 3334 393372 3340
rect 393056 480 393084 3334
rect 394240 3324 394292 3330
rect 394240 3266 394292 3272
rect 394252 480 394280 3266
rect 394712 2774 394740 47670
rect 394804 3602 394832 50102
rect 397012 47734 397040 50102
rect 397472 50102 397854 50130
rect 398852 50102 398958 50130
rect 400062 50102 400168 50130
rect 397000 47728 397052 47734
rect 397000 47670 397052 47676
rect 396540 4140 396592 4146
rect 396540 4082 396592 4088
rect 394792 3596 394844 3602
rect 394792 3538 394844 3544
rect 394712 2746 395384 2774
rect 395356 480 395384 2746
rect 396552 480 396580 4082
rect 397472 3806 397500 50102
rect 398852 45554 398880 50102
rect 400140 47802 400168 50102
rect 400232 50102 401166 50130
rect 401704 50102 402178 50130
rect 403282 50102 403664 50130
rect 404386 50102 404492 50130
rect 405490 50102 405688 50130
rect 406594 50102 406976 50130
rect 400128 47796 400180 47802
rect 400128 47738 400180 47744
rect 399024 47660 399076 47666
rect 399024 47602 399076 47608
rect 398852 45526 398972 45554
rect 398944 16574 398972 45526
rect 398852 16546 398972 16574
rect 398852 4146 398880 16546
rect 398840 4140 398892 4146
rect 398840 4082 398892 4088
rect 397460 3800 397512 3806
rect 397460 3742 397512 3748
rect 397736 3460 397788 3466
rect 397736 3402 397788 3408
rect 397748 480 397776 3402
rect 399036 2774 399064 47602
rect 400232 16574 400260 50102
rect 401600 47864 401652 47870
rect 401600 47806 401652 47812
rect 400232 16546 400352 16574
rect 399116 4140 399168 4146
rect 399116 4082 399168 4088
rect 399128 3942 399156 4082
rect 399116 3936 399168 3942
rect 399116 3878 399168 3884
rect 400128 3868 400180 3874
rect 400128 3810 400180 3816
rect 398944 2746 399064 2774
rect 398944 480 398972 2746
rect 400140 480 400168 3810
rect 400324 3262 400352 16546
rect 401324 3732 401376 3738
rect 401324 3674 401376 3680
rect 400312 3256 400364 3262
rect 400312 3198 400364 3204
rect 401336 480 401364 3674
rect 401612 2774 401640 47806
rect 401704 4146 401732 50102
rect 403636 47666 403664 50102
rect 403624 47660 403676 47666
rect 403624 47602 403676 47608
rect 404464 45554 404492 50102
rect 405660 47870 405688 50102
rect 405648 47864 405700 47870
rect 405648 47806 405700 47812
rect 406948 47598 406976 50102
rect 407132 50102 407698 50130
rect 408604 50102 408802 50130
rect 409800 50102 409906 50130
rect 409984 50102 411010 50130
rect 411272 50102 412114 50130
rect 413218 50102 413600 50130
rect 405740 47592 405792 47598
rect 405740 47534 405792 47540
rect 406936 47592 406988 47598
rect 406936 47534 406988 47540
rect 404372 45526 404492 45554
rect 401692 4140 401744 4146
rect 401692 4082 401744 4088
rect 403624 4004 403676 4010
rect 403624 3946 403676 3952
rect 402980 3664 403032 3670
rect 402980 3606 403032 3612
rect 402992 3330 403020 3606
rect 402980 3324 403032 3330
rect 402980 3266 403032 3272
rect 401612 2746 402560 2774
rect 402532 480 402560 2746
rect 403636 480 403664 3946
rect 404372 3670 404400 45526
rect 405752 16574 405780 47534
rect 405752 16546 406056 16574
rect 404360 3664 404412 3670
rect 404360 3606 404412 3612
rect 404820 3528 404872 3534
rect 404820 3470 404872 3476
rect 404832 480 404860 3470
rect 406028 480 406056 16546
rect 407132 3534 407160 50102
rect 408500 47932 408552 47938
rect 408500 47874 408552 47880
rect 408408 4072 408460 4078
rect 408408 4014 408460 4020
rect 407120 3528 407172 3534
rect 407120 3470 407172 3476
rect 407212 3324 407264 3330
rect 407212 3266 407264 3272
rect 407224 480 407252 3266
rect 408420 480 408448 4014
rect 408512 626 408540 47874
rect 408604 4078 408632 50102
rect 409800 49858 409828 50102
rect 409800 49830 409920 49858
rect 409892 48142 409920 49830
rect 409880 48136 409932 48142
rect 409880 48078 409932 48084
rect 408592 4072 408644 4078
rect 408592 4014 408644 4020
rect 409984 4010 410012 50102
rect 409972 4004 410024 4010
rect 409972 3946 410024 3952
rect 411272 3602 411300 50102
rect 413572 47870 413600 50102
rect 414124 50102 414230 50130
rect 414308 50102 415334 50130
rect 416438 50102 416728 50130
rect 414124 48074 414152 50102
rect 414112 48068 414164 48074
rect 414112 48010 414164 48016
rect 411904 47864 411956 47870
rect 411904 47806 411956 47812
rect 413560 47864 413612 47870
rect 413560 47806 413612 47812
rect 411916 16574 411944 47806
rect 412640 47728 412692 47734
rect 412640 47670 412692 47676
rect 411916 16546 412036 16574
rect 411904 3732 411956 3738
rect 411904 3674 411956 3680
rect 410800 3596 410852 3602
rect 410800 3538 410852 3544
rect 411260 3596 411312 3602
rect 411260 3538 411312 3544
rect 408512 598 409184 626
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 598
rect 410812 480 410840 3538
rect 411916 480 411944 3674
rect 412008 3398 412036 16546
rect 411996 3392 412048 3398
rect 411996 3334 412048 3340
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 47670
rect 414308 45554 414336 50102
rect 416700 48210 416728 50102
rect 416792 50102 417542 50130
rect 418172 50102 418646 50130
rect 419750 50102 420040 50130
rect 416688 48204 416740 48210
rect 416688 48146 416740 48152
rect 415584 47796 415636 47802
rect 415584 47738 415636 47744
rect 414032 45526 414336 45554
rect 414032 3670 414060 45526
rect 415596 16574 415624 47738
rect 415596 16546 416728 16574
rect 415492 3936 415544 3942
rect 415492 3878 415544 3884
rect 414296 3800 414348 3806
rect 414296 3742 414348 3748
rect 414020 3664 414072 3670
rect 414020 3606 414072 3612
rect 414308 480 414336 3742
rect 415504 480 415532 3878
rect 416700 480 416728 16546
rect 416792 3874 416820 50102
rect 416780 3868 416832 3874
rect 416780 3810 416832 3816
rect 418172 3806 418200 50102
rect 420012 48006 420040 50102
rect 420748 50102 420854 50130
rect 420932 50102 421958 50130
rect 423062 50102 423352 50130
rect 420000 48000 420052 48006
rect 420000 47942 420052 47948
rect 420748 47666 420776 50102
rect 419540 47660 419592 47666
rect 419540 47602 419592 47608
rect 420736 47660 420788 47666
rect 420736 47602 420788 47608
rect 419552 16574 419580 47602
rect 419552 16546 420224 16574
rect 418988 4140 419040 4146
rect 418988 4082 419040 4088
rect 418160 3800 418212 3806
rect 418160 3742 418212 3748
rect 417884 3460 417936 3466
rect 417884 3402 417936 3408
rect 417896 480 417924 3402
rect 419000 480 419028 4082
rect 420196 480 420224 16546
rect 420932 3466 420960 50102
rect 423324 47938 423352 50102
rect 423784 50102 424166 50130
rect 425072 50102 425270 50130
rect 426282 50102 426388 50130
rect 427386 50102 427768 50130
rect 423312 47932 423364 47938
rect 423312 47874 423364 47880
rect 423784 16574 423812 50102
rect 423864 47592 423916 47598
rect 423864 47534 423916 47540
rect 423692 16546 423812 16574
rect 423692 3942 423720 16546
rect 423876 6914 423904 47534
rect 423784 6886 423904 6914
rect 423680 3936 423732 3942
rect 423680 3878 423732 3884
rect 421380 3732 421432 3738
rect 421380 3674 421432 3680
rect 420920 3460 420972 3466
rect 420920 3402 420972 3408
rect 421392 480 421420 3674
rect 422576 3392 422628 3398
rect 422576 3334 422628 3340
rect 422588 480 422616 3334
rect 423784 480 423812 6886
rect 425072 3738 425100 50102
rect 426360 47734 426388 50102
rect 426440 48136 426492 48142
rect 426440 48078 426492 48084
rect 426348 47728 426400 47734
rect 426348 47670 426400 47676
rect 426452 16574 426480 48078
rect 427740 47530 427768 50102
rect 427832 50102 428490 50130
rect 429594 50102 429976 50130
rect 430698 50102 430804 50130
rect 427728 47524 427780 47530
rect 427728 47466 427780 47472
rect 426452 16546 426848 16574
rect 426164 4072 426216 4078
rect 426164 4014 426216 4020
rect 425060 3732 425112 3738
rect 425060 3674 425112 3680
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 424980 480 425008 3470
rect 426176 480 426204 4014
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 427832 3534 427860 50102
rect 429948 47598 429976 50102
rect 430580 47864 430632 47870
rect 430776 47818 430804 50102
rect 430580 47806 430632 47812
rect 429936 47592 429988 47598
rect 429936 47534 429988 47540
rect 428464 4004 428516 4010
rect 428464 3946 428516 3952
rect 427820 3528 427872 3534
rect 427820 3470 427872 3476
rect 428476 480 428504 3946
rect 429660 3596 429712 3602
rect 429660 3538 429712 3544
rect 429672 480 429700 3538
rect 430592 3482 430620 47806
rect 430684 47790 430804 47818
rect 431052 50102 431802 50130
rect 432906 50102 433288 50130
rect 434010 50102 434392 50130
rect 430684 3890 430712 47790
rect 431052 45554 431080 50102
rect 433260 48142 433288 50102
rect 434364 48278 434392 50102
rect 434732 50102 435114 50130
rect 436218 50102 436600 50130
rect 437230 50102 437428 50130
rect 438334 50102 438624 50130
rect 439438 50102 439728 50130
rect 434352 48272 434404 48278
rect 434352 48214 434404 48220
rect 433340 48204 433392 48210
rect 433340 48146 433392 48152
rect 433248 48136 433300 48142
rect 433248 48078 433300 48084
rect 432144 48068 432196 48074
rect 432144 48010 432196 48016
rect 430776 45526 431080 45554
rect 430776 4010 430804 45526
rect 432156 6914 432184 48010
rect 433352 16574 433380 48146
rect 433352 16546 434024 16574
rect 432064 6886 432184 6914
rect 430764 4004 430816 4010
rect 430764 3946 430816 3952
rect 430684 3862 430988 3890
rect 430592 3454 430896 3482
rect 430868 480 430896 3454
rect 430960 3398 430988 3862
rect 430948 3392 431000 3398
rect 430948 3334 431000 3340
rect 432064 480 432092 6886
rect 433248 3664 433300 3670
rect 433248 3606 433300 3612
rect 433260 480 433288 3606
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434732 3670 434760 50102
rect 436572 47870 436600 50102
rect 436560 47864 436612 47870
rect 436560 47806 436612 47812
rect 437400 47802 437428 50102
rect 438596 48210 438624 50102
rect 438584 48204 438636 48210
rect 438584 48146 438636 48152
rect 439700 48006 439728 50102
rect 440344 50102 440542 50130
rect 441646 50102 441752 50130
rect 442750 50102 442948 50130
rect 437480 48000 437532 48006
rect 437480 47942 437532 47948
rect 439688 48000 439740 48006
rect 439688 47942 439740 47948
rect 437388 47796 437440 47802
rect 437388 47738 437440 47744
rect 435548 3868 435600 3874
rect 435548 3810 435600 3816
rect 434720 3664 434772 3670
rect 434720 3606 434772 3612
rect 435560 480 435588 3810
rect 436744 3800 436796 3806
rect 436744 3742 436796 3748
rect 436756 480 436784 3742
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 434414 -960 434526 326
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 354 437520 47942
rect 438124 47660 438176 47666
rect 438124 47602 438176 47608
rect 438136 3466 438164 47602
rect 439504 47524 439556 47530
rect 439504 47466 439556 47472
rect 439516 3806 439544 47466
rect 440344 4826 440372 50102
rect 440424 47932 440476 47938
rect 440424 47874 440476 47880
rect 440436 16574 440464 47874
rect 441724 45554 441752 50102
rect 442920 47666 442948 50102
rect 443012 50102 443854 50130
rect 444958 50102 445248 50130
rect 446062 50102 446352 50130
rect 447166 50102 447272 50130
rect 442908 47660 442960 47666
rect 442908 47602 442960 47608
rect 441632 45526 441752 45554
rect 440436 16546 441568 16574
rect 440332 4820 440384 4826
rect 440332 4762 440384 4768
rect 439504 3800 439556 3806
rect 439504 3742 439556 3748
rect 438124 3460 438176 3466
rect 438124 3402 438176 3408
rect 439136 3460 439188 3466
rect 439136 3402 439188 3408
rect 439148 480 439176 3402
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 440344 480 440372 3334
rect 441540 480 441568 16546
rect 441632 4078 441660 45526
rect 441620 4072 441672 4078
rect 441620 4014 441672 4020
rect 442632 3936 442684 3942
rect 442632 3878 442684 3884
rect 442644 480 442672 3878
rect 443012 3602 443040 50102
rect 445220 47938 445248 50102
rect 446324 48074 446352 50102
rect 446404 48272 446456 48278
rect 446404 48214 446456 48220
rect 446312 48068 446364 48074
rect 446312 48010 446364 48016
rect 445208 47932 445260 47938
rect 445208 47874 445260 47880
rect 444380 47728 444432 47734
rect 444380 47670 444432 47676
rect 444392 16574 444420 47670
rect 444392 16546 445064 16574
rect 443828 3732 443880 3738
rect 443828 3674 443880 3680
rect 443000 3596 443052 3602
rect 443000 3538 443052 3544
rect 443840 480 443868 3674
rect 445036 480 445064 16546
rect 446220 3800 446272 3806
rect 446220 3742 446272 3748
rect 446232 480 446260 3742
rect 446416 2990 446444 48214
rect 447244 47818 447272 50102
rect 447152 47790 447272 47818
rect 447428 50102 448270 50130
rect 449282 50102 449664 50130
rect 447152 4146 447180 47790
rect 447428 45554 447456 50102
rect 449636 47734 449664 50102
rect 449912 50102 450386 50130
rect 451490 50102 451872 50130
rect 449624 47728 449676 47734
rect 449624 47670 449676 47676
rect 448612 47592 448664 47598
rect 448612 47534 448664 47540
rect 447244 45526 447456 45554
rect 447140 4140 447192 4146
rect 447140 4082 447192 4088
rect 447244 3942 447272 45526
rect 447232 3936 447284 3942
rect 447232 3878 447284 3884
rect 447416 3528 447468 3534
rect 447416 3470 447468 3476
rect 446404 2984 446456 2990
rect 446404 2926 446456 2932
rect 447428 480 447456 3470
rect 448624 480 448652 47534
rect 449912 3806 449940 50102
rect 451280 48136 451332 48142
rect 451280 48078 451332 48084
rect 451292 16574 451320 48078
rect 451844 47802 451872 50102
rect 452488 50102 452594 50130
rect 452672 50102 453698 50130
rect 454052 50102 454802 50130
rect 455906 50102 456288 50130
rect 457010 50102 457116 50130
rect 451740 47796 451792 47802
rect 451740 47738 451792 47744
rect 451832 47796 451884 47802
rect 451832 47738 451884 47744
rect 451752 47598 451780 47738
rect 451740 47592 451792 47598
rect 451740 47534 451792 47540
rect 452488 47530 452516 50102
rect 452476 47524 452528 47530
rect 452476 47466 452528 47472
rect 451292 16546 451688 16574
rect 450912 4004 450964 4010
rect 450912 3946 450964 3952
rect 449900 3800 449952 3806
rect 449900 3742 449952 3748
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 450924 480 450952 3946
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 452672 3874 452700 50102
rect 453304 47796 453356 47802
rect 453304 47738 453356 47744
rect 452660 3868 452712 3874
rect 452660 3810 452712 3816
rect 453316 3330 453344 47738
rect 454052 3398 454080 50102
rect 454684 48204 454736 48210
rect 454684 48146 454736 48152
rect 454500 3664 454552 3670
rect 454500 3606 454552 3612
rect 454040 3392 454092 3398
rect 454040 3334 454092 3340
rect 453304 3324 453356 3330
rect 453304 3266 453356 3272
rect 453304 2984 453356 2990
rect 453304 2926 453356 2932
rect 453316 480 453344 2926
rect 454512 480 454540 3606
rect 454696 3534 454724 48146
rect 455420 47864 455472 47870
rect 455420 47806 455472 47812
rect 455432 16574 455460 47806
rect 456260 47802 456288 50102
rect 456892 47864 456944 47870
rect 457088 47818 457116 50102
rect 457824 50102 458114 50130
rect 459218 50102 459508 50130
rect 460322 50102 460612 50130
rect 457824 47870 457852 50102
rect 458180 48000 458232 48006
rect 458180 47942 458232 47948
rect 456892 47806 456944 47812
rect 456248 47796 456300 47802
rect 456248 47738 456300 47744
rect 455432 16546 455736 16574
rect 454684 3528 454736 3534
rect 454684 3470 454736 3476
rect 455708 480 455736 16546
rect 456904 6914 456932 47806
rect 456812 6886 456932 6914
rect 456996 47790 457116 47818
rect 457812 47864 457864 47870
rect 457812 47806 457864 47812
rect 456064 4072 456116 4078
rect 456064 4014 456116 4020
rect 456076 3738 456104 4014
rect 456064 3732 456116 3738
rect 456064 3674 456116 3680
rect 456812 3670 456840 6886
rect 456996 4010 457024 47790
rect 457076 47592 457128 47598
rect 457076 47534 457128 47540
rect 456984 4004 457036 4010
rect 456984 3946 457036 3952
rect 456800 3664 456852 3670
rect 456800 3606 456852 3612
rect 457088 3482 457116 47534
rect 458192 16574 458220 47942
rect 459480 47802 459508 50102
rect 460584 48210 460612 50102
rect 460952 50102 461334 50130
rect 462438 50102 462728 50130
rect 463542 50102 463648 50130
rect 460572 48204 460624 48210
rect 460572 48146 460624 48152
rect 459468 47796 459520 47802
rect 459468 47738 459520 47744
rect 458192 16546 459232 16574
rect 458272 3664 458324 3670
rect 458272 3606 458324 3612
rect 456904 3454 457116 3482
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 456904 480 456932 3454
rect 458100 480 458128 3470
rect 458284 3466 458312 3606
rect 458272 3460 458324 3466
rect 458272 3402 458324 3408
rect 459204 480 459232 16546
rect 460388 4820 460440 4826
rect 460388 4762 460440 4768
rect 460400 480 460428 4762
rect 460952 3670 460980 50102
rect 462700 48006 462728 50102
rect 463620 48278 463648 50102
rect 463712 50102 464646 50130
rect 465750 50102 466040 50130
rect 463608 48272 463660 48278
rect 463608 48214 463660 48220
rect 462688 48000 462740 48006
rect 462688 47942 462740 47948
rect 462320 47660 462372 47666
rect 462320 47602 462372 47608
rect 461584 3732 461636 3738
rect 461584 3674 461636 3680
rect 460940 3664 460992 3670
rect 460940 3606 460992 3612
rect 461596 480 461624 3674
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 354 462360 47602
rect 463712 3738 463740 50102
rect 465264 48068 465316 48074
rect 465264 48010 465316 48016
rect 464344 47932 464396 47938
rect 464344 47874 464396 47880
rect 463700 3732 463752 3738
rect 463700 3674 463752 3680
rect 464356 3602 464384 47874
rect 465276 16574 465304 48010
rect 466012 47938 466040 50102
rect 466472 50102 466854 50130
rect 467958 50102 468248 50130
rect 469062 50102 469168 50130
rect 466000 47932 466052 47938
rect 466000 47874 466052 47880
rect 465276 16546 465856 16574
rect 463976 3596 464028 3602
rect 463976 3538 464028 3544
rect 464344 3596 464396 3602
rect 464344 3538 464396 3544
rect 465172 3596 465224 3602
rect 465172 3538 465224 3544
rect 463988 480 464016 3538
rect 465184 480 465212 3538
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 466472 4962 466500 50102
rect 468220 47666 468248 50102
rect 469140 48142 469168 50102
rect 469324 50102 470166 50130
rect 470612 50102 471270 50130
rect 472282 50102 472664 50130
rect 473386 50102 473492 50130
rect 474490 50102 474688 50130
rect 475594 50102 475976 50130
rect 469128 48136 469180 48142
rect 469128 48078 469180 48084
rect 469220 47728 469272 47734
rect 469220 47670 469272 47676
rect 468208 47660 468260 47666
rect 468208 47602 468260 47608
rect 466460 4956 466512 4962
rect 466460 4898 466512 4904
rect 467472 4140 467524 4146
rect 467472 4082 467524 4088
rect 467484 480 467512 4082
rect 468668 3936 468720 3942
rect 468668 3878 468720 3884
rect 468680 480 468708 3878
rect 469232 3482 469260 47670
rect 469324 5166 469352 50102
rect 469312 5160 469364 5166
rect 469312 5102 469364 5108
rect 470612 3602 470640 50102
rect 472636 47734 472664 50102
rect 472624 47728 472676 47734
rect 472624 47670 472676 47676
rect 473464 16574 473492 50102
rect 474660 48074 474688 50102
rect 474648 48068 474700 48074
rect 474648 48010 474700 48016
rect 475384 47864 475436 47870
rect 475384 47806 475436 47812
rect 473544 47592 473596 47598
rect 473544 47534 473596 47540
rect 473372 16546 473492 16574
rect 473372 5234 473400 16546
rect 473556 6914 473584 47534
rect 473464 6886 473584 6914
rect 473360 5228 473412 5234
rect 473360 5170 473412 5176
rect 471060 3800 471112 3806
rect 471060 3742 471112 3748
rect 470600 3596 470652 3602
rect 470600 3538 470652 3544
rect 469232 3454 469904 3482
rect 469876 480 469904 3454
rect 471072 480 471100 3742
rect 472256 3392 472308 3398
rect 472256 3334 472308 3340
rect 472268 480 472296 3334
rect 473464 480 473492 6886
rect 474556 3868 474608 3874
rect 474556 3810 474608 3816
rect 474568 480 474596 3810
rect 475396 3534 475424 47806
rect 475948 47598 475976 50102
rect 476132 50102 476698 50130
rect 477802 50102 478184 50130
rect 478906 50102 479012 50130
rect 475936 47592 475988 47598
rect 475936 47534 475988 47540
rect 476132 4894 476160 50102
rect 478052 48272 478104 48278
rect 478052 48214 478104 48220
rect 476764 48204 476816 48210
rect 476764 48146 476816 48152
rect 476120 4888 476172 4894
rect 476120 4830 476172 4836
rect 475384 3528 475436 3534
rect 475384 3470 475436 3476
rect 475752 3460 475804 3466
rect 475752 3402 475804 3408
rect 475764 480 475792 3402
rect 476776 3058 476804 48146
rect 478064 45554 478092 48214
rect 478156 48210 478184 50102
rect 478144 48204 478196 48210
rect 478144 48146 478196 48152
rect 478984 47784 479012 50102
rect 478892 47756 479012 47784
rect 479076 50102 480010 50130
rect 481114 50102 481496 50130
rect 482218 50102 482600 50130
rect 478064 45526 478184 45554
rect 478156 16574 478184 45526
rect 478156 16546 478276 16574
rect 478144 4004 478196 4010
rect 478144 3946 478196 3952
rect 476948 3528 477000 3534
rect 476948 3470 477000 3476
rect 476764 3052 476816 3058
rect 476764 2994 476816 3000
rect 476960 480 476988 3470
rect 478156 480 478184 3946
rect 478248 3534 478276 16546
rect 478892 5030 478920 47756
rect 479076 45554 479104 50102
rect 481272 47932 481324 47938
rect 481272 47874 481324 47880
rect 480260 47796 480312 47802
rect 480260 47738 480312 47744
rect 478984 45526 479104 45554
rect 478880 5024 478932 5030
rect 478880 4966 478932 4972
rect 478984 4826 479012 45526
rect 480272 16574 480300 47738
rect 481284 47530 481312 47874
rect 481468 47870 481496 50102
rect 482284 48068 482336 48074
rect 482284 48010 482336 48016
rect 481456 47864 481508 47870
rect 481456 47806 481508 47812
rect 481272 47524 481324 47530
rect 481272 47466 481324 47472
rect 480272 16546 480576 16574
rect 478972 4820 479024 4826
rect 478972 4762 479024 4768
rect 478236 3528 478288 3534
rect 478236 3470 478288 3476
rect 479340 3392 479392 3398
rect 479340 3334 479392 3340
rect 479352 480 479380 3334
rect 480548 480 480576 16546
rect 482296 3806 482324 48010
rect 482572 47938 482600 50102
rect 483216 50102 483322 50130
rect 483400 50102 484334 50130
rect 485438 50102 485728 50130
rect 483020 48068 483072 48074
rect 483020 48010 483072 48016
rect 482560 47932 482612 47938
rect 482560 47874 482612 47880
rect 482284 3800 482336 3806
rect 482284 3742 482336 3748
rect 482836 3664 482888 3670
rect 482836 3606 482888 3612
rect 481732 3052 481784 3058
rect 481732 2994 481784 3000
rect 481744 480 481772 2994
rect 482848 480 482876 3606
rect 483032 3482 483060 48010
rect 483216 48006 483244 50102
rect 483204 48000 483256 48006
rect 483204 47942 483256 47948
rect 483400 45554 483428 50102
rect 485044 48204 485096 48210
rect 485044 48146 485096 48152
rect 483124 45526 483428 45554
rect 483124 3670 483152 45526
rect 485056 4146 485084 48146
rect 485700 47802 485728 50102
rect 485792 50102 486542 50130
rect 487646 50102 487936 50130
rect 485688 47796 485740 47802
rect 485688 47738 485740 47744
rect 485044 4140 485096 4146
rect 485044 4082 485096 4088
rect 483112 3664 483164 3670
rect 483112 3606 483164 3612
rect 485792 3534 485820 50102
rect 486424 47864 486476 47870
rect 486424 47806 486476 47812
rect 486436 3942 486464 47806
rect 487160 47524 487212 47530
rect 487160 47466 487212 47472
rect 486424 3936 486476 3942
rect 486424 3878 486476 3884
rect 486424 3732 486476 3738
rect 486424 3674 486476 3680
rect 485228 3528 485280 3534
rect 483032 3454 484072 3482
rect 485228 3470 485280 3476
rect 485780 3528 485832 3534
rect 485780 3470 485832 3476
rect 484044 480 484072 3454
rect 485240 480 485268 3470
rect 486436 480 486464 3674
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 47466
rect 487908 46986 487936 50102
rect 488644 50102 488750 50130
rect 488828 50102 489854 50130
rect 490116 50102 490958 50130
rect 492062 50102 492352 50130
rect 488644 48074 488672 50102
rect 488632 48068 488684 48074
rect 488632 48010 488684 48016
rect 487896 46980 487948 46986
rect 487896 46922 487948 46928
rect 488828 45554 488856 50102
rect 489920 48136 489972 48142
rect 489920 48078 489972 48084
rect 488552 45526 488856 45554
rect 488552 5098 488580 45526
rect 488540 5092 488592 5098
rect 488540 5034 488592 5040
rect 488816 4956 488868 4962
rect 488816 4898 488868 4904
rect 488828 480 488856 4898
rect 489932 3466 489960 48078
rect 490012 47660 490064 47666
rect 490012 47602 490064 47608
rect 489920 3460 489972 3466
rect 489920 3402 489972 3408
rect 490024 3346 490052 47602
rect 490116 3398 490144 50102
rect 492324 47938 492352 50102
rect 492692 50102 493166 50130
rect 494270 50102 494560 50130
rect 492312 47932 492364 47938
rect 492312 47874 492364 47880
rect 490564 46980 490616 46986
rect 490564 46922 490616 46928
rect 490576 4078 490604 46922
rect 492312 5160 492364 5166
rect 492312 5102 492364 5108
rect 490564 4072 490616 4078
rect 490564 4014 490616 4020
rect 490748 3460 490800 3466
rect 490748 3402 490800 3408
rect 489932 3318 490052 3346
rect 490104 3392 490156 3398
rect 490104 3334 490156 3340
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3402
rect 492324 480 492352 5102
rect 492692 4010 492720 50102
rect 494532 48142 494560 50102
rect 495268 50102 495374 50130
rect 495452 50102 496386 50130
rect 496832 50102 497490 50130
rect 498594 50102 498976 50130
rect 494520 48136 494572 48142
rect 494520 48078 494572 48084
rect 495268 47734 495296 50102
rect 494060 47728 494112 47734
rect 494060 47670 494112 47676
rect 495256 47728 495308 47734
rect 495256 47670 495308 47676
rect 494072 16574 494100 47670
rect 494072 16546 494744 16574
rect 492680 4004 492732 4010
rect 492680 3946 492732 3952
rect 493508 3596 493560 3602
rect 493508 3538 493560 3544
rect 493520 480 493548 3538
rect 494716 480 494744 16546
rect 495452 4962 495480 50102
rect 495900 5228 495952 5234
rect 495900 5170 495952 5176
rect 495440 4956 495492 4962
rect 495440 4898 495492 4904
rect 495912 480 495940 5170
rect 496832 3602 496860 50102
rect 498948 47666 498976 50102
rect 499592 50102 499698 50130
rect 499776 50102 500802 50130
rect 501906 50102 502288 50130
rect 498936 47660 498988 47666
rect 498936 47602 498988 47608
rect 498200 47592 498252 47598
rect 498200 47534 498252 47540
rect 497096 3800 497148 3806
rect 497096 3742 497148 3748
rect 496820 3596 496872 3602
rect 496820 3538 496872 3544
rect 497108 480 497136 3742
rect 498212 480 498240 47534
rect 499396 4888 499448 4894
rect 499396 4830 499448 4836
rect 499408 480 499436 4830
rect 499592 3874 499620 50102
rect 499580 3868 499632 3874
rect 499580 3810 499632 3816
rect 499776 3806 499804 50102
rect 502260 47598 502288 50102
rect 502352 50102 503010 50130
rect 503732 50102 504114 50130
rect 505218 50102 505324 50130
rect 502248 47592 502300 47598
rect 502248 47534 502300 47540
rect 502352 5030 502380 50102
rect 501788 5024 501840 5030
rect 501788 4966 501840 4972
rect 502340 5024 502392 5030
rect 502340 4966 502392 4972
rect 500592 4140 500644 4146
rect 500592 4082 500644 4088
rect 499764 3800 499816 3806
rect 499764 3742 499816 3748
rect 500604 480 500632 4082
rect 501800 480 501828 4966
rect 502984 4820 503036 4826
rect 502984 4762 503036 4768
rect 502996 480 503024 4762
rect 503732 3738 503760 50102
rect 505100 47864 505152 47870
rect 505296 47818 505324 50102
rect 505100 47806 505152 47812
rect 504180 3936 504232 3942
rect 504180 3878 504232 3884
rect 503720 3732 503772 3738
rect 503720 3674 503772 3680
rect 504192 480 504220 3878
rect 505112 3482 505140 47806
rect 505204 47790 505324 47818
rect 505388 50102 506322 50130
rect 506584 50102 507426 50130
rect 508438 50102 508728 50130
rect 505204 5234 505232 47790
rect 505388 45554 505416 50102
rect 505296 45526 505416 45554
rect 505192 5228 505244 5234
rect 505192 5170 505244 5176
rect 505296 4894 505324 45526
rect 505284 4888 505336 4894
rect 505284 4830 505336 4836
rect 506584 3942 506612 50102
rect 508700 48006 508728 50102
rect 509252 50102 509542 50130
rect 510646 50102 510752 50130
rect 506664 48000 506716 48006
rect 506664 47942 506716 47948
rect 508688 48000 508740 48006
rect 508688 47942 508740 47948
rect 506572 3936 506624 3942
rect 506572 3878 506624 3884
rect 505112 3454 505416 3482
rect 505388 480 505416 3454
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 354 506562 480
rect 506676 354 506704 47942
rect 507860 47796 507912 47802
rect 507860 47738 507912 47744
rect 507872 16574 507900 47738
rect 507872 16546 508912 16574
rect 507676 3664 507728 3670
rect 507676 3606 507728 3612
rect 507688 480 507716 3606
rect 508884 480 508912 16546
rect 509252 5166 509280 50102
rect 510724 47818 510752 50102
rect 510632 47790 510752 47818
rect 510816 50102 511750 50130
rect 512104 50102 512854 50130
rect 513958 50102 514248 50130
rect 515062 50102 515352 50130
rect 516166 50102 516272 50130
rect 517270 50102 517468 50130
rect 509240 5160 509292 5166
rect 509240 5102 509292 5108
rect 510632 3670 510660 47790
rect 510816 45554 510844 50102
rect 512000 48068 512052 48074
rect 512000 48010 512052 48016
rect 510724 45526 510844 45554
rect 510724 4826 510752 45526
rect 510712 4820 510764 4826
rect 510712 4762 510764 4768
rect 511264 4072 511316 4078
rect 511264 4014 511316 4020
rect 510620 3664 510672 3670
rect 510620 3606 510672 3612
rect 510068 3528 510120 3534
rect 510068 3470 510120 3476
rect 510080 480 510108 3470
rect 511276 480 511304 4014
rect 506450 326 506704 354
rect 506450 -960 506562 326
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 48010
rect 512104 3534 512132 50102
rect 514220 48210 514248 50102
rect 514208 48204 514260 48210
rect 514208 48146 514260 48152
rect 515324 48074 515352 50102
rect 515404 48136 515456 48142
rect 515404 48078 515456 48084
rect 515312 48068 515364 48074
rect 515312 48010 515364 48016
rect 514852 47932 514904 47938
rect 514852 47874 514904 47880
rect 514864 16574 514892 47874
rect 514864 16546 515352 16574
rect 513564 5092 513616 5098
rect 513564 5034 513616 5040
rect 512092 3528 512144 3534
rect 512092 3470 512144 3476
rect 513576 480 513604 5034
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515324 490 515352 16546
rect 515416 3058 515444 48078
rect 516244 45554 516272 50102
rect 517440 47938 517468 50102
rect 517532 50102 518374 50130
rect 519386 50102 519768 50130
rect 517428 47932 517480 47938
rect 517428 47874 517480 47880
rect 516152 45526 516272 45554
rect 516152 5506 516180 45526
rect 516140 5500 516192 5506
rect 516140 5442 516192 5448
rect 517532 5370 517560 50102
rect 518900 47728 518952 47734
rect 518900 47670 518952 47676
rect 518912 16574 518940 47670
rect 519740 47394 519768 50102
rect 520292 50102 520490 50130
rect 521488 50102 521594 50130
rect 522698 50102 522988 50130
rect 519728 47388 519780 47394
rect 519728 47330 519780 47336
rect 518912 16546 519584 16574
rect 517520 5364 517572 5370
rect 517520 5306 517572 5312
rect 517152 4004 517204 4010
rect 517152 3946 517204 3952
rect 515404 3052 515456 3058
rect 515404 2994 515456 3000
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515324 462 515536 490
rect 517164 480 517192 3946
rect 518348 3052 518400 3058
rect 518348 2994 518400 3000
rect 518360 480 518388 2994
rect 519556 480 519584 16546
rect 520292 3466 520320 50102
rect 521488 47530 521516 50102
rect 521476 47524 521528 47530
rect 521476 47466 521528 47472
rect 522304 47388 522356 47394
rect 522304 47330 522356 47336
rect 520740 4956 520792 4962
rect 520740 4898 520792 4904
rect 520280 3460 520332 3466
rect 520280 3402 520332 3408
rect 520752 480 520780 4898
rect 522316 4010 522344 47330
rect 522960 47326 522988 50102
rect 523144 50102 523802 50130
rect 524906 50102 525288 50130
rect 526010 50102 526116 50130
rect 522948 47320 523000 47326
rect 522948 47262 523000 47268
rect 523144 4146 523172 50102
rect 525064 48204 525116 48210
rect 525064 48146 525116 48152
rect 523224 47660 523276 47666
rect 523224 47602 523276 47608
rect 523132 4140 523184 4146
rect 523132 4082 523184 4088
rect 522304 4004 522356 4010
rect 522304 3946 522356 3952
rect 521844 3596 521896 3602
rect 521844 3538 521896 3544
rect 521856 480 521884 3538
rect 515508 354 515536 462
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 354 523122 480
rect 523236 354 523264 47602
rect 524328 4140 524380 4146
rect 524328 4082 524380 4088
rect 524340 3874 524368 4082
rect 524236 3868 524288 3874
rect 524236 3810 524288 3816
rect 524328 3868 524380 3874
rect 524328 3810 524380 3816
rect 524248 480 524276 3810
rect 525076 3602 525104 48146
rect 525260 47802 525288 50102
rect 525892 47864 525944 47870
rect 525892 47806 525944 47812
rect 525248 47796 525300 47802
rect 525248 47738 525300 47744
rect 525800 47592 525852 47598
rect 525800 47534 525852 47540
rect 525432 3800 525484 3806
rect 525432 3742 525484 3748
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 525444 480 525472 3742
rect 525812 490 525840 47534
rect 525904 3806 525932 47806
rect 526088 45554 526116 50102
rect 526824 50102 527114 50130
rect 528218 50102 528324 50130
rect 526824 47870 526852 50102
rect 526812 47864 526864 47870
rect 526812 47806 526864 47812
rect 528296 47666 528324 50102
rect 528572 50102 529322 50130
rect 530426 50102 530808 50130
rect 528284 47660 528336 47666
rect 528284 47602 528336 47608
rect 525996 45526 526116 45554
rect 525996 5438 526024 45526
rect 525984 5432 526036 5438
rect 525984 5374 526036 5380
rect 528572 5098 528600 50102
rect 530780 48142 530808 50102
rect 531332 50102 531438 50130
rect 531516 50102 532542 50130
rect 532804 50102 533646 50130
rect 534750 50102 535040 50130
rect 535854 50102 536144 50130
rect 536958 50102 537248 50130
rect 530768 48136 530820 48142
rect 530768 48078 530820 48084
rect 529204 47320 529256 47326
rect 529204 47262 529256 47268
rect 528560 5092 528612 5098
rect 528560 5034 528612 5040
rect 527824 5024 527876 5030
rect 527824 4966 527876 4972
rect 525892 3800 525944 3806
rect 525892 3742 525944 3748
rect 523010 326 523264 354
rect 523010 -960 523122 326
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 525812 462 526208 490
rect 527836 480 527864 4966
rect 529216 4078 529244 47262
rect 531332 5302 531360 50102
rect 531320 5296 531372 5302
rect 531320 5238 531372 5244
rect 531516 5234 531544 50102
rect 532700 48000 532752 48006
rect 532700 47942 532752 47948
rect 530124 5228 530176 5234
rect 530124 5170 530176 5176
rect 531504 5228 531556 5234
rect 531504 5170 531556 5176
rect 529204 4072 529256 4078
rect 529204 4014 529256 4020
rect 529020 3732 529072 3738
rect 529020 3674 529072 3680
rect 529032 480 529060 3674
rect 530136 480 530164 5170
rect 531320 4888 531372 4894
rect 531320 4830 531372 4836
rect 531332 480 531360 4830
rect 532516 3936 532568 3942
rect 532516 3878 532568 3884
rect 532528 480 532556 3878
rect 532712 3482 532740 47942
rect 532804 3738 532832 50102
rect 535012 47598 535040 50102
rect 536116 47734 536144 50102
rect 537220 48006 537248 50102
rect 537588 50102 538062 50130
rect 538232 50102 539166 50130
rect 539704 50102 540270 50130
rect 540992 50102 541374 50130
rect 542478 50102 542584 50130
rect 543490 50102 543688 50130
rect 537208 48000 537260 48006
rect 537208 47942 537260 47948
rect 536104 47728 536156 47734
rect 536104 47670 536156 47676
rect 535000 47592 535052 47598
rect 535000 47534 535052 47540
rect 537588 45554 537616 50102
rect 536852 45526 537616 45554
rect 534908 5160 534960 5166
rect 534908 5102 534960 5108
rect 532792 3732 532844 3738
rect 532792 3674 532844 3680
rect 532712 3454 533752 3482
rect 533724 480 533752 3454
rect 534920 480 534948 5102
rect 536852 4962 536880 45526
rect 538232 5030 538260 50102
rect 538220 5024 538272 5030
rect 538220 4966 538272 4972
rect 536840 4956 536892 4962
rect 536840 4898 536892 4904
rect 537208 4820 537260 4826
rect 537208 4762 537260 4768
rect 536104 3664 536156 3670
rect 536104 3606 536156 3612
rect 536116 480 536144 3606
rect 537220 480 537248 4762
rect 539704 3670 539732 50102
rect 539784 48068 539836 48074
rect 539784 48010 539836 48016
rect 539796 16574 539824 48010
rect 539796 16546 540376 16574
rect 539692 3664 539744 3670
rect 539692 3606 539744 3612
rect 539600 3596 539652 3602
rect 539600 3538 539652 3544
rect 538404 3528 538456 3534
rect 538404 3470 538456 3476
rect 538416 480 538444 3470
rect 539612 480 539640 3538
rect 526180 354 526208 462
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 540992 4894 541020 50102
rect 542360 47932 542412 47938
rect 542360 47874 542412 47880
rect 541992 5500 542044 5506
rect 541992 5442 542044 5448
rect 540980 4888 541032 4894
rect 540980 4830 541032 4836
rect 542004 480 542032 5442
rect 542372 490 542400 47874
rect 542556 45554 542584 50102
rect 543660 47938 543688 50102
rect 543752 50102 544594 50130
rect 545132 50102 545698 50130
rect 546512 50102 546802 50130
rect 547906 50102 548288 50130
rect 549010 50102 549208 50130
rect 550114 50102 550496 50130
rect 551218 50102 551600 50130
rect 552322 50102 552704 50130
rect 553426 50102 553532 50130
rect 543648 47932 543700 47938
rect 543648 47874 543700 47880
rect 542464 45526 542584 45554
rect 542464 5166 542492 45526
rect 542452 5160 542504 5166
rect 542452 5102 542504 5108
rect 543752 4826 543780 50102
rect 544384 5364 544436 5370
rect 544384 5306 544436 5312
rect 543740 4820 543792 4826
rect 543740 4762 543792 4768
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542372 462 542768 490
rect 544396 480 544424 5306
rect 545132 3534 545160 50102
rect 545488 4004 545540 4010
rect 545488 3946 545540 3952
rect 545120 3528 545172 3534
rect 545120 3470 545172 3476
rect 545500 480 545528 3946
rect 546512 3602 546540 50102
rect 548260 47938 548288 50102
rect 548156 47932 548208 47938
rect 548156 47874 548208 47880
rect 548248 47932 548300 47938
rect 548248 47874 548300 47880
rect 548168 47530 548196 47874
rect 549180 47870 549208 50102
rect 550468 48006 550496 50102
rect 550456 48000 550508 48006
rect 550456 47942 550508 47948
rect 549168 47864 549220 47870
rect 549168 47806 549220 47812
rect 551284 47864 551336 47870
rect 551284 47806 551336 47812
rect 550640 47796 550692 47802
rect 550640 47738 550692 47744
rect 548064 47524 548116 47530
rect 548064 47466 548116 47472
rect 548156 47524 548208 47530
rect 548156 47466 548208 47472
rect 546500 3596 546552 3602
rect 546500 3538 546552 3544
rect 546684 3460 546736 3466
rect 546684 3402 546736 3408
rect 546696 480 546724 3402
rect 542740 354 542768 462
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 354 547962 480
rect 548076 354 548104 47466
rect 550652 16574 550680 47738
rect 550652 16546 551048 16574
rect 549076 4072 549128 4078
rect 549076 4014 549128 4020
rect 549088 480 549116 4014
rect 550272 3868 550324 3874
rect 550272 3810 550324 3816
rect 550284 480 550312 3810
rect 547850 326 548104 354
rect 547850 -960 547962 326
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 551296 3874 551324 47806
rect 551572 47394 551600 50102
rect 552676 47870 552704 50102
rect 552664 47864 552716 47870
rect 552664 47806 552716 47812
rect 551560 47388 551612 47394
rect 551560 47330 551612 47336
rect 553504 45554 553532 50102
rect 554044 48136 554096 48142
rect 554044 48078 554096 48084
rect 553412 45526 553532 45554
rect 552664 5432 552716 5438
rect 552664 5374 552716 5380
rect 551284 3868 551336 3874
rect 551284 3810 551336 3816
rect 552676 480 552704 5374
rect 553412 3466 553440 45526
rect 553768 3800 553820 3806
rect 553768 3742 553820 3748
rect 553400 3460 553452 3466
rect 553400 3402 553452 3408
rect 553780 480 553808 3742
rect 554056 3194 554084 48078
rect 555424 48068 555476 48074
rect 555424 48010 555476 48016
rect 554780 47660 554832 47666
rect 554780 47602 554832 47608
rect 554044 3188 554096 3194
rect 554044 3130 554096 3136
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 47602
rect 555436 4146 555464 48010
rect 556896 48000 556948 48006
rect 556896 47942 556948 47948
rect 556804 47524 556856 47530
rect 556804 47466 556856 47472
rect 556160 5092 556212 5098
rect 556160 5034 556212 5040
rect 555424 4140 555476 4146
rect 555424 4082 555476 4088
rect 556172 480 556200 5034
rect 556816 4078 556844 47466
rect 556804 4072 556856 4078
rect 556804 4014 556856 4020
rect 556908 3942 556936 47942
rect 560944 47864 560996 47870
rect 560944 47806 560996 47812
rect 558184 47388 558236 47394
rect 558184 47330 558236 47336
rect 556896 3936 556948 3942
rect 556896 3878 556948 3884
rect 558196 3806 558224 47330
rect 558552 5296 558604 5302
rect 558552 5238 558604 5244
rect 558184 3800 558236 3806
rect 558184 3742 558236 3748
rect 557356 3188 557408 3194
rect 557356 3130 557408 3136
rect 557368 480 557396 3130
rect 558564 480 558592 5238
rect 559748 5228 559800 5234
rect 559748 5170 559800 5176
rect 559760 480 559788 5170
rect 560956 4010 560984 47806
rect 566464 47796 566516 47802
rect 566464 47738 566516 47744
rect 563060 47728 563112 47734
rect 563060 47670 563112 47676
rect 561680 47592 561732 47598
rect 561680 47534 561732 47540
rect 561692 16574 561720 47534
rect 561692 16546 562088 16574
rect 560944 4004 560996 4010
rect 560944 3946 560996 3952
rect 560852 3732 560904 3738
rect 560852 3674 560904 3680
rect 560864 480 560892 3674
rect 562060 480 562088 16546
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 47670
rect 565636 4956 565688 4962
rect 565636 4898 565688 4904
rect 564440 4140 564492 4146
rect 564440 4082 564492 4088
rect 564452 480 564480 4082
rect 565648 480 565676 4898
rect 566476 3738 566504 47738
rect 570328 5160 570380 5166
rect 570328 5102 570380 5108
rect 566832 5024 566884 5030
rect 566832 4966 566884 4972
rect 566464 3732 566516 3738
rect 566464 3674 566516 3680
rect 566844 480 566872 4966
rect 569132 4888 569184 4894
rect 569132 4830 569184 4836
rect 568028 3664 568080 3670
rect 568028 3606 568080 3612
rect 568040 480 568068 3606
rect 569144 480 569172 4830
rect 570340 480 570368 5102
rect 572720 4820 572772 4826
rect 572720 4762 572772 4768
rect 571524 4072 571576 4078
rect 571524 4014 571576 4020
rect 571536 480 571564 4014
rect 572732 480 572760 4762
rect 582196 4004 582248 4010
rect 582196 3946 582248 3952
rect 578608 3936 578660 3942
rect 578608 3878 578660 3884
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 576308 3732 576360 3738
rect 576308 3674 576360 3680
rect 575112 3596 575164 3602
rect 575112 3538 575164 3544
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 573928 480 573956 3470
rect 575124 480 575152 3538
rect 576320 480 576348 3674
rect 577424 480 577452 3810
rect 578620 480 578648 3878
rect 581000 3800 581052 3806
rect 581000 3742 581052 3748
rect 581012 480 581040 3742
rect 582208 480 582236 3946
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3698 673784 3754 673840
rect 3606 673648 3662 673704
rect 3238 671200 3294 671256
rect 3146 658180 3148 658200
rect 3148 658180 3200 658200
rect 3200 658180 3202 658200
rect 3146 658144 3202 658180
rect 3146 632032 3202 632088
rect 3238 619112 3294 619168
rect 3146 606056 3202 606112
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3330 553832 3386 553888
rect 3238 501744 3294 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 3146 449556 3148 449576
rect 3148 449556 3200 449576
rect 3200 449556 3202 449576
rect 3146 449520 3202 449556
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3146 397432 3202 397488
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 2778 345344 2834 345400
rect 2778 306212 2780 306232
rect 2780 306212 2832 306232
rect 2832 306212 2834 306232
rect 2778 306176 2834 306212
rect 2778 254088 2834 254144
rect 2778 201864 2834 201920
rect 4802 672560 4858 672616
rect 4066 514800 4122 514856
rect 3974 319232 4030 319288
rect 3882 293120 3938 293176
rect 3790 267144 3846 267200
rect 3698 241032 3754 241088
rect 3606 214920 3662 214976
rect 3514 188808 3570 188864
rect 3422 162832 3478 162888
rect 2778 149776 2834 149832
rect 3238 136720 3294 136776
rect 2778 97552 2834 97608
rect 2778 84632 2834 84688
rect 4986 672288 5042 672344
rect 6458 668072 6514 668128
rect 11702 673512 11758 673568
rect 44822 670792 44878 670848
rect 68190 672424 68246 672480
rect 101126 673920 101182 673976
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 471426 673784 471482 673840
rect 397090 672424 397146 672480
rect 396354 671064 396410 671120
rect 438950 670928 439006 670984
rect 448150 669976 448206 670032
rect 485778 673648 485834 673704
rect 499578 673512 499634 673568
rect 532698 672560 532754 672616
rect 518346 672288 518402 672344
rect 523130 671200 523186 671256
rect 139490 669568 139546 669624
rect 162122 669568 162178 669624
rect 358910 669568 358966 669624
rect 35438 669432 35494 669488
rect 16486 669296 16542 669352
rect 21270 669296 21326 669352
rect 25962 669296 26018 669352
rect 30654 669296 30710 669352
rect 39946 669296 40002 669352
rect 527730 669296 527786 669352
rect 537114 669296 537170 669352
rect 541898 669296 541954 669352
rect 546590 669296 546646 669352
rect 556802 673920 556858 673976
rect 579618 670656 579674 670712
rect 580078 668480 580134 668536
rect 579986 644000 580042 644056
rect 579986 630808 580042 630864
rect 579986 617480 580042 617536
rect 579802 590960 579858 591016
rect 579802 577632 579858 577688
rect 579986 564340 579988 564360
rect 579988 564340 580040 564360
rect 580040 564340 580042 564360
rect 579986 564304 580042 564340
rect 579986 537784 580042 537840
rect 579986 524456 580042 524512
rect 579986 511264 580042 511320
rect 579802 471416 579858 471472
rect 579986 458124 579988 458144
rect 579988 458124 580040 458144
rect 580040 458124 580042 458144
rect 579986 458088 580042 458124
rect 579986 431568 580042 431624
rect 579986 418240 580042 418296
rect 579986 404912 580042 404968
rect 579802 378392 579858 378448
rect 579986 365064 580042 365120
rect 579986 351872 580042 351928
rect 579986 325216 580042 325272
rect 579986 312024 580042 312080
rect 580078 298696 580134 298752
rect 580078 272176 580134 272232
rect 580078 258848 580134 258904
rect 580078 245556 580080 245576
rect 580080 245556 580132 245576
rect 580132 245556 580134 245576
rect 580078 245520 580134 245556
rect 580262 669296 580318 669352
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 579618 165824 579674 165880
rect 579618 125976 579674 126032
rect 580906 205672 580962 205728
rect 580814 192480 580870 192536
rect 580722 179152 580778 179208
rect 580630 152632 580686 152688
rect 580538 139304 580594 139360
rect 580446 112784 580502 112840
rect 580354 99456 580410 99512
rect 580262 59608 580318 59664
rect 2778 58520 2834 58576
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 101121 673978 101187 673981
rect 556797 673978 556863 673981
rect 101121 673976 556863 673978
rect 101121 673920 101126 673976
rect 101182 673920 556802 673976
rect 556858 673920 556863 673976
rect 101121 673918 556863 673920
rect 101121 673915 101187 673918
rect 556797 673915 556863 673918
rect 3693 673842 3759 673845
rect 471421 673842 471487 673845
rect 3693 673840 471487 673842
rect 3693 673784 3698 673840
rect 3754 673784 471426 673840
rect 471482 673784 471487 673840
rect 3693 673782 471487 673784
rect 3693 673779 3759 673782
rect 471421 673779 471487 673782
rect 3601 673706 3667 673709
rect 485773 673706 485839 673709
rect 3601 673704 485839 673706
rect 3601 673648 3606 673704
rect 3662 673648 485778 673704
rect 485834 673648 485839 673704
rect 3601 673646 485839 673648
rect 3601 673643 3667 673646
rect 485773 673643 485839 673646
rect 11697 673570 11763 673573
rect 499573 673570 499639 673573
rect 11697 673568 499639 673570
rect 11697 673512 11702 673568
rect 11758 673512 499578 673568
rect 499634 673512 499639 673568
rect 11697 673510 499639 673512
rect 11697 673507 11763 673510
rect 499573 673507 499639 673510
rect 4797 672618 4863 672621
rect 532693 672618 532759 672621
rect 4797 672616 532759 672618
rect 4797 672560 4802 672616
rect 4858 672560 532698 672616
rect 532754 672560 532759 672616
rect 4797 672558 532759 672560
rect 4797 672555 4863 672558
rect 532693 672555 532759 672558
rect 68185 672482 68251 672485
rect 397085 672482 397151 672485
rect 68185 672480 397151 672482
rect 68185 672424 68190 672480
rect 68246 672424 397090 672480
rect 397146 672424 397151 672480
rect 68185 672422 397151 672424
rect 68185 672419 68251 672422
rect 397085 672419 397151 672422
rect 4981 672346 5047 672349
rect 518341 672346 518407 672349
rect 4981 672344 518407 672346
rect 4981 672288 4986 672344
rect 5042 672288 518346 672344
rect 518402 672288 518407 672344
rect 4981 672286 518407 672288
rect 4981 672283 5047 672286
rect 518341 672283 518407 672286
rect -960 671258 480 671348
rect 3233 671258 3299 671261
rect 523125 671258 523191 671261
rect -960 671256 3299 671258
rect -960 671200 3238 671256
rect 3294 671200 3299 671256
rect -960 671198 3299 671200
rect -960 671108 480 671198
rect 3233 671195 3299 671198
rect 6870 671256 523191 671258
rect 6870 671200 523130 671256
rect 523186 671200 523191 671256
rect 6870 671198 523191 671200
rect 3366 671060 3372 671124
rect 3436 671122 3442 671124
rect 6870 671122 6930 671198
rect 523125 671195 523191 671198
rect 3436 671062 6930 671122
rect 3436 671060 3442 671062
rect 14590 671060 14596 671124
rect 14660 671122 14666 671124
rect 396349 671122 396415 671125
rect 14660 671120 396415 671122
rect 14660 671064 396354 671120
rect 396410 671064 396415 671120
rect 14660 671062 396415 671064
rect 14660 671060 14666 671062
rect 396349 671059 396415 671062
rect 14406 670924 14412 670988
rect 14476 670986 14482 670988
rect 438945 670986 439011 670989
rect 14476 670984 439011 670986
rect 14476 670928 438950 670984
rect 439006 670928 439011 670984
rect 14476 670926 439011 670928
rect 14476 670924 14482 670926
rect 438945 670923 439011 670926
rect 44817 670850 44883 670853
rect 554078 670850 554084 670852
rect 44817 670848 554084 670850
rect 44817 670792 44822 670848
rect 44878 670792 554084 670848
rect 44817 670790 554084 670792
rect 44817 670787 44883 670790
rect 554078 670788 554084 670790
rect 554148 670788 554154 670852
rect 579613 670714 579679 670717
rect 583520 670714 584960 670804
rect 579613 670712 584960 670714
rect 579613 670656 579618 670712
rect 579674 670656 584960 670712
rect 579613 670654 584960 670656
rect 579613 670651 579679 670654
rect 583520 670564 584960 670654
rect 448145 670034 448211 670037
rect 431910 670032 448211 670034
rect 431910 669976 448150 670032
rect 448206 669976 448211 670032
rect 431910 669974 448211 669976
rect 3550 669836 3556 669900
rect 3620 669898 3626 669900
rect 431910 669898 431970 669974
rect 448145 669971 448211 669974
rect 3620 669838 431970 669898
rect 3620 669836 3626 669838
rect 139485 669628 139551 669629
rect 162117 669628 162183 669629
rect 358905 669628 358971 669629
rect 139485 669626 139532 669628
rect 139440 669624 139532 669626
rect 139440 669568 139490 669624
rect 139440 669566 139532 669568
rect 139485 669564 139532 669566
rect 139596 669564 139602 669628
rect 162117 669624 162164 669628
rect 162228 669626 162234 669628
rect 358854 669626 358860 669628
rect 162117 669568 162122 669624
rect 162117 669564 162164 669568
rect 162228 669566 162274 669626
rect 358814 669566 358860 669626
rect 358924 669624 358971 669628
rect 358966 669568 358971 669624
rect 162228 669564 162234 669566
rect 358854 669564 358860 669566
rect 358924 669564 358971 669568
rect 139485 669563 139551 669564
rect 162117 669563 162183 669564
rect 358905 669563 358971 669564
rect 35433 669490 35499 669493
rect 553894 669490 553900 669492
rect 35433 669488 553900 669490
rect 35433 669432 35438 669488
rect 35494 669432 553900 669488
rect 35433 669430 553900 669432
rect 35433 669427 35499 669430
rect 553894 669428 553900 669430
rect 553964 669428 553970 669492
rect 16481 669356 16547 669357
rect 16430 669354 16436 669356
rect 16390 669294 16436 669354
rect 16500 669352 16547 669356
rect 16542 669296 16547 669352
rect 16430 669292 16436 669294
rect 16500 669292 16547 669296
rect 16481 669291 16547 669292
rect 21265 669354 21331 669357
rect 25957 669356 26023 669357
rect 21950 669354 21956 669356
rect 21265 669352 21956 669354
rect 21265 669296 21270 669352
rect 21326 669296 21956 669352
rect 21265 669294 21956 669296
rect 21265 669291 21331 669294
rect 21950 669292 21956 669294
rect 22020 669292 22026 669356
rect 25957 669352 26004 669356
rect 26068 669354 26074 669356
rect 30649 669354 30715 669357
rect 30782 669354 30788 669356
rect 25957 669296 25962 669352
rect 25957 669292 26004 669296
rect 26068 669294 26114 669354
rect 30649 669352 30788 669354
rect 30649 669296 30654 669352
rect 30710 669296 30788 669352
rect 30649 669294 30788 669296
rect 26068 669292 26074 669294
rect 25957 669291 26023 669292
rect 30649 669291 30715 669294
rect 30782 669292 30788 669294
rect 30852 669292 30858 669356
rect 39941 669354 40007 669357
rect 39941 669352 527098 669354
rect 39941 669296 39946 669352
rect 40002 669296 527098 669352
rect 39941 669294 527098 669296
rect 39941 669291 40007 669294
rect 527038 669218 527098 669294
rect 527214 669292 527220 669356
rect 527284 669354 527290 669356
rect 527725 669354 527791 669357
rect 527284 669352 527791 669354
rect 527284 669296 527730 669352
rect 527786 669296 527791 669352
rect 527284 669294 527791 669296
rect 527284 669292 527290 669294
rect 527725 669291 527791 669294
rect 527958 669294 536666 669354
rect 527958 669218 528018 669294
rect 527038 669158 528018 669218
rect 536606 669218 536666 669294
rect 536782 669292 536788 669356
rect 536852 669354 536858 669356
rect 537109 669354 537175 669357
rect 536852 669352 537175 669354
rect 536852 669296 537114 669352
rect 537170 669296 537175 669352
rect 536852 669294 537175 669296
rect 536852 669292 536858 669294
rect 537109 669291 537175 669294
rect 537342 669294 540898 669354
rect 537342 669218 537402 669294
rect 536606 669158 537402 669218
rect 540838 669218 540898 669294
rect 541014 669292 541020 669356
rect 541084 669354 541090 669356
rect 541893 669354 541959 669357
rect 546585 669356 546651 669357
rect 546534 669354 546540 669356
rect 541084 669352 541959 669354
rect 541084 669296 541898 669352
rect 541954 669296 541959 669352
rect 541084 669294 541959 669296
rect 541084 669292 541090 669294
rect 541893 669291 541959 669294
rect 542126 669294 546418 669354
rect 546494 669294 546540 669354
rect 546604 669352 546651 669356
rect 580257 669354 580323 669357
rect 546646 669296 546651 669352
rect 542126 669218 542186 669294
rect 540838 669158 542186 669218
rect 546358 669218 546418 669294
rect 546534 669292 546540 669294
rect 546604 669292 546651 669296
rect 546585 669291 546651 669292
rect 546726 669352 580323 669354
rect 546726 669296 580262 669352
rect 580318 669296 580323 669352
rect 546726 669294 580323 669296
rect 546726 669218 546786 669294
rect 580257 669291 580323 669294
rect 546358 669158 546786 669218
rect 139526 668476 139532 668540
rect 139596 668538 139602 668540
rect 580073 668538 580139 668541
rect 139596 668536 580139 668538
rect 139596 668480 580078 668536
rect 580134 668480 580139 668536
rect 139596 668478 580139 668480
rect 139596 668476 139602 668478
rect 580073 668475 580139 668478
rect 6453 668130 6519 668133
rect 358854 668130 358860 668132
rect 6453 668128 358860 668130
rect 6453 668072 6458 668128
rect 6514 668072 358860 668128
rect 6453 668070 358860 668072
rect 6453 668067 6519 668070
rect 358854 668068 358860 668070
rect 358924 668068 358930 668132
rect 162158 667932 162164 667996
rect 162228 667994 162234 667996
rect 540094 667994 540100 667996
rect 162228 667934 540100 667994
rect 162228 667932 162234 667934
rect 540094 667932 540100 667934
rect 540164 667932 540170 667996
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 579981 644058 580047 644061
rect 583520 644058 584960 644148
rect 579981 644056 584960 644058
rect 579981 644000 579986 644056
rect 580042 644000 584960 644056
rect 579981 643998 584960 644000
rect 579981 643995 580047 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3141 632090 3207 632093
rect -960 632088 3207 632090
rect -960 632032 3146 632088
rect 3202 632032 3207 632088
rect -960 632030 3207 632032
rect -960 631940 480 632030
rect 3141 632027 3207 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3233 619170 3299 619173
rect -960 619168 3299 619170
rect -960 619112 3238 619168
rect 3294 619112 3299 619168
rect -960 619110 3299 619112
rect -960 619020 480 619110
rect 3233 619107 3299 619110
rect 579981 617538 580047 617541
rect 583520 617538 584960 617628
rect 579981 617536 584960 617538
rect 579981 617480 579986 617536
rect 580042 617480 584960 617536
rect 579981 617478 584960 617480
rect 579981 617475 580047 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3141 606114 3207 606117
rect -960 606112 3207 606114
rect -960 606056 3146 606112
rect 3202 606056 3207 606112
rect -960 606054 3207 606056
rect -960 605964 480 606054
rect 3141 606051 3207 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 579797 577690 579863 577693
rect 583520 577690 584960 577780
rect 579797 577688 584960 577690
rect 579797 577632 579802 577688
rect 579858 577632 584960 577688
rect 579797 577630 584960 577632
rect 579797 577627 579863 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 579981 564362 580047 564365
rect 583520 564362 584960 564452
rect 579981 564360 584960 564362
rect 579981 564304 579986 564360
rect 580042 564304 584960 564360
rect 579981 564302 584960 564304
rect 579981 564299 580047 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579981 537842 580047 537845
rect 583520 537842 584960 537932
rect 579981 537840 584960 537842
rect 579981 537784 579986 537840
rect 580042 537784 584960 537840
rect 579981 537782 584960 537784
rect 579981 537779 580047 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect -960 527854 674 527914
rect -960 527778 480 527854
rect 614 527778 674 527854
rect -960 527764 674 527778
rect 246 527718 674 527764
rect 246 527234 306 527718
rect 13854 527234 13860 527236
rect 246 527174 13860 527234
rect 13854 527172 13860 527174
rect 13924 527172 13930 527236
rect 579981 524514 580047 524517
rect 583520 524514 584960 524604
rect 579981 524512 584960 524514
rect 579981 524456 579986 524512
rect 580042 524456 584960 524512
rect 579981 524454 584960 524456
rect 579981 524451 580047 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 4061 514858 4127 514861
rect -960 514856 4127 514858
rect -960 514800 4066 514856
rect 4122 514800 4127 514856
rect -960 514798 4127 514800
rect -960 514708 480 514798
rect 4061 514795 4127 514798
rect 579981 511322 580047 511325
rect 583520 511322 584960 511412
rect 579981 511320 584960 511322
rect 579981 511264 579986 511320
rect 580042 511264 584960 511320
rect 579981 511262 584960 511264
rect 579981 511259 580047 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484666 584960 484756
rect 567150 484606 584960 484666
rect 541014 484468 541020 484532
rect 541084 484530 541090 484532
rect 567150 484530 567210 484606
rect 541084 484470 567210 484530
rect 583520 484516 584960 484606
rect 541084 484468 541090 484470
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 579797 471474 579863 471477
rect 583520 471474 584960 471564
rect 579797 471472 584960 471474
rect 579797 471416 579802 471472
rect 579858 471416 584960 471472
rect 579797 471414 584960 471416
rect 579797 471411 579863 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 579981 458146 580047 458149
rect 583520 458146 584960 458236
rect 579981 458144 584960 458146
rect 579981 458088 579986 458144
rect 580042 458088 584960 458144
rect 579981 458086 584960 458088
rect 579981 458083 580047 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579981 431626 580047 431629
rect 583520 431626 584960 431716
rect 579981 431624 584960 431626
rect 579981 431568 579986 431624
rect 580042 431568 584960 431624
rect 579981 431566 584960 431568
rect 579981 431563 580047 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579981 418298 580047 418301
rect 583520 418298 584960 418388
rect 579981 418296 584960 418298
rect 579981 418240 579986 418296
rect 580042 418240 584960 418296
rect 579981 418238 584960 418240
rect 579981 418235 580047 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3141 397490 3207 397493
rect -960 397488 3207 397490
rect -960 397432 3146 397488
rect 3202 397432 3207 397488
rect -960 397430 3207 397432
rect -960 397340 480 397430
rect 3141 397427 3207 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 13854 371378 13860 371380
rect -960 371318 13860 371378
rect -960 371228 480 371318
rect 13854 371316 13860 371318
rect 13924 371316 13930 371380
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 579981 365059 580047 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 579981 351930 580047 351933
rect 583520 351930 584960 352020
rect 579981 351928 584960 351930
rect 579981 351872 579986 351928
rect 580042 351872 584960 351928
rect 579981 351870 584960 351872
rect 579981 351867 580047 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3969 319290 4035 319293
rect -960 319288 4035 319290
rect -960 319232 3974 319288
rect 4030 319232 4035 319288
rect -960 319230 4035 319232
rect -960 319140 480 319230
rect 3969 319227 4035 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 2773 306234 2839 306237
rect -960 306232 2839 306234
rect -960 306176 2778 306232
rect 2834 306176 2839 306232
rect -960 306174 2839 306176
rect -960 306084 480 306174
rect 2773 306171 2839 306174
rect 580073 298754 580139 298757
rect 583520 298754 584960 298844
rect 580073 298752 584960 298754
rect 580073 298696 580078 298752
rect 580134 298696 584960 298752
rect 580073 298694 584960 298696
rect 580073 298691 580139 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3877 293178 3943 293181
rect -960 293176 3943 293178
rect -960 293120 3882 293176
rect 3938 293120 3943 293176
rect -960 293118 3943 293120
rect -960 293028 480 293118
rect 3877 293115 3943 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580073 272234 580139 272237
rect 583520 272234 584960 272324
rect 580073 272232 584960 272234
rect 580073 272176 580078 272232
rect 580134 272176 584960 272232
rect 580073 272174 584960 272176
rect 580073 272171 580139 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3785 267202 3851 267205
rect -960 267200 3851 267202
rect -960 267144 3790 267200
rect 3846 267144 3851 267200
rect -960 267142 3851 267144
rect -960 267052 480 267142
rect 3785 267139 3851 267142
rect 580073 258906 580139 258909
rect 583520 258906 584960 258996
rect 580073 258904 584960 258906
rect 580073 258848 580078 258904
rect 580134 258848 584960 258904
rect 580073 258846 584960 258848
rect 580073 258843 580139 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 580073 245578 580139 245581
rect 583520 245578 584960 245668
rect 580073 245576 584960 245578
rect 580073 245520 580078 245576
rect 580134 245520 584960 245576
rect 580073 245518 584960 245520
rect 580073 245515 580139 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3693 241090 3759 241093
rect -960 241088 3759 241090
rect -960 241032 3698 241088
rect 3754 241032 3759 241088
rect -960 241030 3759 241032
rect -960 240940 480 241030
rect 3693 241027 3759 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3601 214978 3667 214981
rect -960 214976 3667 214978
rect -960 214920 3606 214976
rect 3662 214920 3667 214976
rect -960 214918 3667 214920
rect -960 214828 480 214918
rect 3601 214915 3667 214918
rect 580901 205730 580967 205733
rect 583520 205730 584960 205820
rect 580901 205728 584960 205730
rect 580901 205672 580906 205728
rect 580962 205672 584960 205728
rect 580901 205670 584960 205672
rect 580901 205667 580967 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580809 192538 580875 192541
rect 583520 192538 584960 192628
rect 580809 192536 584960 192538
rect 580809 192480 580814 192536
rect 580870 192480 584960 192536
rect 580809 192478 584960 192480
rect 580809 192475 580875 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 580717 179210 580783 179213
rect 583520 179210 584960 179300
rect 580717 179208 584960 179210
rect 580717 179152 580722 179208
rect 580778 179152 584960 179208
rect 580717 179150 584960 179152
rect 580717 179147 580783 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 579613 165882 579679 165885
rect 583520 165882 584960 165972
rect 579613 165880 584960 165882
rect 579613 165824 579618 165880
rect 579674 165824 584960 165880
rect 579613 165822 584960 165824
rect 579613 165819 579679 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 580625 152690 580691 152693
rect 583520 152690 584960 152780
rect 580625 152688 584960 152690
rect 580625 152632 580630 152688
rect 580686 152632 584960 152688
rect 580625 152630 584960 152632
rect 580625 152627 580691 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 580533 139362 580599 139365
rect 583520 139362 584960 139452
rect 580533 139360 584960 139362
rect 580533 139304 580538 139360
rect 580594 139304 584960 139360
rect 580533 139302 584960 139304
rect 580533 139299 580599 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3550 110666 3556 110668
rect -960 110606 3556 110666
rect -960 110516 480 110606
rect 3550 110604 3556 110606
rect 3620 110604 3626 110668
rect 580349 99514 580415 99517
rect 583520 99514 584960 99604
rect 580349 99512 584960 99514
rect 580349 99456 580354 99512
rect 580410 99456 584960 99512
rect 580349 99454 584960 99456
rect 580349 99451 580415 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 554078 85580 554084 85644
rect 554148 85642 554154 85644
rect 583526 85642 583586 85990
rect 554148 85582 583586 85642
rect 554148 85580 554154 85582
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 553894 71844 553900 71908
rect 553964 71906 553970 71908
rect 583526 71906 583586 72798
rect 553964 71846 583586 71906
rect 553964 71844 553970 71846
rect -960 71634 480 71724
rect 3366 71634 3372 71636
rect -960 71574 3372 71634
rect -960 71484 480 71574
rect 3366 71572 3372 71574
rect 3436 71572 3442 71636
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2773 58578 2839 58581
rect -960 58576 2839 58578
rect -960 58520 2778 58576
rect 2834 58520 2839 58576
rect -960 58518 2839 58520
rect -960 58428 480 58518
rect 2773 58515 2839 58518
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect -960 45522 480 45612
rect 30782 45596 30788 45660
rect 30852 45658 30858 45660
rect 583526 45658 583586 46142
rect 30852 45598 583586 45658
rect 30852 45596 30858 45598
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 527214 44298 527220 44300
rect 6870 44238 527220 44298
rect 527214 44236 527220 44238
rect 527284 44236 527290 44300
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31922 306 32270
rect 536782 31922 536788 31924
rect 246 31862 536788 31922
rect 536782 31860 536788 31862
rect 536852 31860 536858 31924
rect 21950 31724 21956 31788
rect 22020 31786 22026 31788
rect 583526 31786 583586 32950
rect 22020 31726 583586 31786
rect 22020 31724 22026 31726
rect 583520 19818 584960 19908
rect 583342 19758 584960 19818
rect 583342 19682 583402 19758
rect 583520 19682 584960 19758
rect 583342 19668 584960 19682
rect 583342 19622 583586 19668
rect 546534 19546 546540 19548
rect -960 19410 480 19500
rect 6870 19486 546540 19546
rect 6870 19410 6930 19486
rect 546534 19484 546540 19486
rect 546604 19484 546610 19548
rect -960 19350 6930 19410
rect -960 19260 480 19350
rect 25998 19348 26004 19412
rect 26068 19410 26074 19412
rect 583526 19410 583586 19622
rect 26068 19350 583586 19410
rect 26068 19348 26074 19350
rect 583520 6626 584960 6716
rect -960 6490 480 6580
rect 583342 6566 584960 6626
rect 583342 6490 583402 6566
rect 583520 6490 584960 6566
rect -960 6430 674 6490
rect 583342 6476 584960 6490
rect 583342 6430 583586 6476
rect -960 6354 480 6430
rect 614 6354 674 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 246 5810 306 6294
rect 541014 5810 541020 5812
rect 246 5750 541020 5810
rect 541014 5748 541020 5750
rect 541084 5748 541090 5812
rect 16430 5612 16436 5676
rect 16500 5674 16506 5676
rect 583526 5674 583586 6430
rect 16500 5614 583586 5674
rect 16500 5612 16506 5614
<< via3 >>
rect 3372 671060 3436 671124
rect 14596 671060 14660 671124
rect 14412 670924 14476 670988
rect 554084 670788 554148 670852
rect 3556 669836 3620 669900
rect 139532 669624 139596 669628
rect 139532 669568 139546 669624
rect 139546 669568 139596 669624
rect 139532 669564 139596 669568
rect 162164 669624 162228 669628
rect 162164 669568 162178 669624
rect 162178 669568 162228 669624
rect 162164 669564 162228 669568
rect 358860 669624 358924 669628
rect 358860 669568 358910 669624
rect 358910 669568 358924 669624
rect 358860 669564 358924 669568
rect 553900 669428 553964 669492
rect 16436 669352 16500 669356
rect 16436 669296 16486 669352
rect 16486 669296 16500 669352
rect 16436 669292 16500 669296
rect 21956 669292 22020 669356
rect 26004 669352 26068 669356
rect 26004 669296 26018 669352
rect 26018 669296 26068 669352
rect 26004 669292 26068 669296
rect 30788 669292 30852 669356
rect 527220 669292 527284 669356
rect 536788 669292 536852 669356
rect 541020 669292 541084 669356
rect 546540 669352 546604 669356
rect 546540 669296 546590 669352
rect 546590 669296 546604 669352
rect 546540 669292 546604 669296
rect 139532 668476 139596 668540
rect 358860 668068 358924 668132
rect 162164 667932 162228 667996
rect 540100 667932 540164 667996
rect 13860 527172 13924 527236
rect 541020 484468 541084 484532
rect 13860 371316 13924 371380
rect 3556 110604 3620 110668
rect 554084 85580 554148 85644
rect 553900 71844 553964 71908
rect 3372 71572 3436 71636
rect 30788 45596 30852 45660
rect 527220 44236 527284 44300
rect 536788 31860 536852 31924
rect 21956 31724 22020 31788
rect 546540 19484 546604 19548
rect 26004 19348 26068 19412
rect 541020 5748 541084 5812
rect 16436 5612 16500 5676
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3371 671124 3437 671125
rect 3371 671060 3372 671124
rect 3436 671060 3437 671124
rect 3371 671059 3437 671060
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 71637 3434 671059
rect 3555 669900 3621 669901
rect 3555 669836 3556 669900
rect 3620 669836 3621 669900
rect 3555 669835 3621 669836
rect 3558 110669 3618 669835
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3555 110668 3621 110669
rect 3555 110604 3556 110668
rect 3620 110604 3621 110668
rect 3555 110603 3621 110604
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3371 71636 3437 71637
rect 3371 71572 3372 71636
rect 3436 71572 3437 71636
rect 3371 71571 3437 71572
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 672000 13574 698058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 672000 20414 705242
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 672000 24134 672618
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 672000 27854 676338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 672000 31574 680058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 672000 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 672000 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 672000 45854 694338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 672000 49574 698058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 672000 56414 705242
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 672000 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 672000 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 672000 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 672000 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 672000 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 672000 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 672000 85574 698058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 672000 92414 705242
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 672000 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 672000 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 672000 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 672000 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 672000 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 672000 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 672000 121574 698058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 672000 128414 705242
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 672000 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 672000 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 672000 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 672000 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 672000 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 672000 153854 694338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 672000 157574 698058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 672000 164414 705242
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 672000 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 672000 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 672000 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 672000 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 672000 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 672000 189854 694338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 672000 193574 698058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 672000 200414 705242
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 672000 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 672000 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 672000 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 672000 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 672000 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 672000 225854 694338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 672000 229574 698058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 672000 236414 705242
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 672000 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 672000 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 672000 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 672000 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 672000 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 672000 261854 694338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 672000 265574 698058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 672000 272414 705242
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 672000 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 672000 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 672000 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 672000 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 672000 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 672000 297854 694338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 672000 301574 698058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 672000 308414 705242
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 672000 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 672000 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 672000 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 672000 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 672000 330134 690618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 672000 333854 694338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 672000 337574 698058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 672000 344414 705242
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 672000 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 672000 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 672000 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 672000 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 672000 366134 690618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 672000 369854 694338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 672000 373574 698058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 672000 380414 705242
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 672000 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 672000 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 672000 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 672000 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 672000 402134 690618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 672000 405854 694338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 672000 409574 698058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 672000 416414 705242
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 672000 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 672000 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 672000 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 672000 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 672000 438134 690618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 672000 441854 694338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 672000 445574 698058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 672000 452414 705242
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 672000 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 672000 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 672000 463574 680058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 672000 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 672000 474134 690618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 672000 477854 694338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 672000 481574 698058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 672000 488414 705242
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 672000 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 672000 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 672000 499574 680058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 672000 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 672000 510134 690618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 672000 513854 694338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 672000 517574 698058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 672000 524414 705242
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 672000 528134 672618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 672000 531854 676338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 672000 535574 680058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 672000 542414 686898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 672000 546134 690618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 672000 549854 694338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 672000 553574 698058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 14595 671124 14661 671125
rect 14595 671060 14596 671124
rect 14660 671060 14661 671124
rect 14595 671059 14661 671060
rect 14411 670988 14477 670989
rect 14411 670924 14412 670988
rect 14476 670924 14477 670988
rect 14411 670923 14477 670924
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 14414 534090 14474 670923
rect 14230 534030 14474 534090
rect 14230 531330 14290 534030
rect 13678 531270 14290 531330
rect 13678 521670 13738 531270
rect 13859 527236 13925 527237
rect 13859 527172 13860 527236
rect 13924 527234 13925 527236
rect 14598 527234 14658 671059
rect 554083 670852 554149 670853
rect 554083 670788 554084 670852
rect 554148 670788 554149 670852
rect 554083 670787 554149 670788
rect 139531 669628 139597 669629
rect 139531 669564 139532 669628
rect 139596 669564 139597 669628
rect 139531 669563 139597 669564
rect 162163 669628 162229 669629
rect 162163 669564 162164 669628
rect 162228 669564 162229 669628
rect 162163 669563 162229 669564
rect 358859 669628 358925 669629
rect 358859 669564 358860 669628
rect 358924 669564 358925 669628
rect 358859 669563 358925 669564
rect 16435 669356 16501 669357
rect 16435 669292 16436 669356
rect 16500 669292 16501 669356
rect 16435 669291 16501 669292
rect 21955 669356 22021 669357
rect 21955 669292 21956 669356
rect 22020 669292 22021 669356
rect 21955 669291 22021 669292
rect 26003 669356 26069 669357
rect 26003 669292 26004 669356
rect 26068 669292 26069 669356
rect 26003 669291 26069 669292
rect 30787 669356 30853 669357
rect 30787 669292 30788 669356
rect 30852 669292 30853 669356
rect 30787 669291 30853 669292
rect 13924 527174 14658 527234
rect 13924 527172 13925 527174
rect 13859 527171 13925 527172
rect 13678 521610 14474 521670
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 14414 374010 14474 521610
rect 13862 373950 14474 374010
rect 13862 371381 13922 373950
rect 13859 371380 13925 371381
rect 13859 371316 13860 371380
rect 13924 371316 13925 371380
rect 13859 371315 13925 371316
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 14614 13574 48000
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 16438 5677 16498 669291
rect 18208 651454 18528 651486
rect 18208 651218 18250 651454
rect 18486 651218 18528 651454
rect 18208 651134 18528 651218
rect 18208 650898 18250 651134
rect 18486 650898 18528 651134
rect 18208 650866 18528 650898
rect 18208 615454 18528 615486
rect 18208 615218 18250 615454
rect 18486 615218 18528 615454
rect 18208 615134 18528 615218
rect 18208 614898 18250 615134
rect 18486 614898 18528 615134
rect 18208 614866 18528 614898
rect 18208 579454 18528 579486
rect 18208 579218 18250 579454
rect 18486 579218 18528 579454
rect 18208 579134 18528 579218
rect 18208 578898 18250 579134
rect 18486 578898 18528 579134
rect 18208 578866 18528 578898
rect 18208 543454 18528 543486
rect 18208 543218 18250 543454
rect 18486 543218 18528 543454
rect 18208 543134 18528 543218
rect 18208 542898 18250 543134
rect 18486 542898 18528 543134
rect 18208 542866 18528 542898
rect 18208 507454 18528 507486
rect 18208 507218 18250 507454
rect 18486 507218 18528 507454
rect 18208 507134 18528 507218
rect 18208 506898 18250 507134
rect 18486 506898 18528 507134
rect 18208 506866 18528 506898
rect 18208 471454 18528 471486
rect 18208 471218 18250 471454
rect 18486 471218 18528 471454
rect 18208 471134 18528 471218
rect 18208 470898 18250 471134
rect 18486 470898 18528 471134
rect 18208 470866 18528 470898
rect 18208 435454 18528 435486
rect 18208 435218 18250 435454
rect 18486 435218 18528 435454
rect 18208 435134 18528 435218
rect 18208 434898 18250 435134
rect 18486 434898 18528 435134
rect 18208 434866 18528 434898
rect 18208 399454 18528 399486
rect 18208 399218 18250 399454
rect 18486 399218 18528 399454
rect 18208 399134 18528 399218
rect 18208 398898 18250 399134
rect 18486 398898 18528 399134
rect 18208 398866 18528 398898
rect 18208 363454 18528 363486
rect 18208 363218 18250 363454
rect 18486 363218 18528 363454
rect 18208 363134 18528 363218
rect 18208 362898 18250 363134
rect 18486 362898 18528 363134
rect 18208 362866 18528 362898
rect 18208 327454 18528 327486
rect 18208 327218 18250 327454
rect 18486 327218 18528 327454
rect 18208 327134 18528 327218
rect 18208 326898 18250 327134
rect 18486 326898 18528 327134
rect 18208 326866 18528 326898
rect 18208 291454 18528 291486
rect 18208 291218 18250 291454
rect 18486 291218 18528 291454
rect 18208 291134 18528 291218
rect 18208 290898 18250 291134
rect 18486 290898 18528 291134
rect 18208 290866 18528 290898
rect 18208 255454 18528 255486
rect 18208 255218 18250 255454
rect 18486 255218 18528 255454
rect 18208 255134 18528 255218
rect 18208 254898 18250 255134
rect 18486 254898 18528 255134
rect 18208 254866 18528 254898
rect 18208 219454 18528 219486
rect 18208 219218 18250 219454
rect 18486 219218 18528 219454
rect 18208 219134 18528 219218
rect 18208 218898 18250 219134
rect 18486 218898 18528 219134
rect 18208 218866 18528 218898
rect 18208 183454 18528 183486
rect 18208 183218 18250 183454
rect 18486 183218 18528 183454
rect 18208 183134 18528 183218
rect 18208 182898 18250 183134
rect 18486 182898 18528 183134
rect 18208 182866 18528 182898
rect 18208 147454 18528 147486
rect 18208 147218 18250 147454
rect 18486 147218 18528 147454
rect 18208 147134 18528 147218
rect 18208 146898 18250 147134
rect 18486 146898 18528 147134
rect 18208 146866 18528 146898
rect 18208 111454 18528 111486
rect 18208 111218 18250 111454
rect 18486 111218 18528 111454
rect 18208 111134 18528 111218
rect 18208 110898 18250 111134
rect 18486 110898 18528 111134
rect 18208 110866 18528 110898
rect 18208 75454 18528 75486
rect 18208 75218 18250 75454
rect 18486 75218 18528 75454
rect 18208 75134 18528 75218
rect 18208 74898 18250 75134
rect 18486 74898 18528 75134
rect 18208 74866 18528 74898
rect 19794 21454 20414 48000
rect 21958 31789 22018 669291
rect 21955 31788 22021 31789
rect 21955 31724 21956 31788
rect 22020 31724 22021 31788
rect 21955 31723 22021 31724
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 16435 5676 16501 5677
rect 16435 5612 16436 5676
rect 16500 5612 16501 5676
rect 16435 5611 16501 5612
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 25174 24134 48000
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 26006 19413 26066 669291
rect 27234 28894 27854 48000
rect 30790 45661 30850 669291
rect 139534 668541 139594 669563
rect 139531 668540 139597 668541
rect 139531 668476 139532 668540
rect 139596 668476 139597 668540
rect 139531 668475 139597 668476
rect 162166 667997 162226 669563
rect 358862 668133 358922 669563
rect 553899 669492 553965 669493
rect 553899 669428 553900 669492
rect 553964 669428 553965 669492
rect 553899 669427 553965 669428
rect 527219 669356 527285 669357
rect 527219 669292 527220 669356
rect 527284 669292 527285 669356
rect 527219 669291 527285 669292
rect 536787 669356 536853 669357
rect 536787 669292 536788 669356
rect 536852 669292 536853 669356
rect 536787 669291 536853 669292
rect 541019 669356 541085 669357
rect 541019 669292 541020 669356
rect 541084 669292 541085 669356
rect 541019 669291 541085 669292
rect 546539 669356 546605 669357
rect 546539 669292 546540 669356
rect 546604 669292 546605 669356
rect 546539 669291 546605 669292
rect 358859 668132 358925 668133
rect 358859 668068 358860 668132
rect 358924 668068 358925 668132
rect 358859 668067 358925 668068
rect 162163 667996 162229 667997
rect 162163 667932 162164 667996
rect 162228 667932 162229 667996
rect 162163 667931 162229 667932
rect 48928 651454 49248 651486
rect 48928 651218 48970 651454
rect 49206 651218 49248 651454
rect 48928 651134 49248 651218
rect 48928 650898 48970 651134
rect 49206 650898 49248 651134
rect 48928 650866 49248 650898
rect 79648 651454 79968 651486
rect 79648 651218 79690 651454
rect 79926 651218 79968 651454
rect 79648 651134 79968 651218
rect 79648 650898 79690 651134
rect 79926 650898 79968 651134
rect 79648 650866 79968 650898
rect 110368 651454 110688 651486
rect 110368 651218 110410 651454
rect 110646 651218 110688 651454
rect 110368 651134 110688 651218
rect 110368 650898 110410 651134
rect 110646 650898 110688 651134
rect 110368 650866 110688 650898
rect 141088 651454 141408 651486
rect 141088 651218 141130 651454
rect 141366 651218 141408 651454
rect 141088 651134 141408 651218
rect 141088 650898 141130 651134
rect 141366 650898 141408 651134
rect 141088 650866 141408 650898
rect 171808 651454 172128 651486
rect 171808 651218 171850 651454
rect 172086 651218 172128 651454
rect 171808 651134 172128 651218
rect 171808 650898 171850 651134
rect 172086 650898 172128 651134
rect 171808 650866 172128 650898
rect 202528 651454 202848 651486
rect 202528 651218 202570 651454
rect 202806 651218 202848 651454
rect 202528 651134 202848 651218
rect 202528 650898 202570 651134
rect 202806 650898 202848 651134
rect 202528 650866 202848 650898
rect 233248 651454 233568 651486
rect 233248 651218 233290 651454
rect 233526 651218 233568 651454
rect 233248 651134 233568 651218
rect 233248 650898 233290 651134
rect 233526 650898 233568 651134
rect 233248 650866 233568 650898
rect 263968 651454 264288 651486
rect 263968 651218 264010 651454
rect 264246 651218 264288 651454
rect 263968 651134 264288 651218
rect 263968 650898 264010 651134
rect 264246 650898 264288 651134
rect 263968 650866 264288 650898
rect 294688 651454 295008 651486
rect 294688 651218 294730 651454
rect 294966 651218 295008 651454
rect 294688 651134 295008 651218
rect 294688 650898 294730 651134
rect 294966 650898 295008 651134
rect 294688 650866 295008 650898
rect 325408 651454 325728 651486
rect 325408 651218 325450 651454
rect 325686 651218 325728 651454
rect 325408 651134 325728 651218
rect 325408 650898 325450 651134
rect 325686 650898 325728 651134
rect 325408 650866 325728 650898
rect 356128 651454 356448 651486
rect 356128 651218 356170 651454
rect 356406 651218 356448 651454
rect 356128 651134 356448 651218
rect 356128 650898 356170 651134
rect 356406 650898 356448 651134
rect 356128 650866 356448 650898
rect 386848 651454 387168 651486
rect 386848 651218 386890 651454
rect 387126 651218 387168 651454
rect 386848 651134 387168 651218
rect 386848 650898 386890 651134
rect 387126 650898 387168 651134
rect 386848 650866 387168 650898
rect 417568 651454 417888 651486
rect 417568 651218 417610 651454
rect 417846 651218 417888 651454
rect 417568 651134 417888 651218
rect 417568 650898 417610 651134
rect 417846 650898 417888 651134
rect 417568 650866 417888 650898
rect 448288 651454 448608 651486
rect 448288 651218 448330 651454
rect 448566 651218 448608 651454
rect 448288 651134 448608 651218
rect 448288 650898 448330 651134
rect 448566 650898 448608 651134
rect 448288 650866 448608 650898
rect 479008 651454 479328 651486
rect 479008 651218 479050 651454
rect 479286 651218 479328 651454
rect 479008 651134 479328 651218
rect 479008 650898 479050 651134
rect 479286 650898 479328 651134
rect 479008 650866 479328 650898
rect 509728 651454 510048 651486
rect 509728 651218 509770 651454
rect 510006 651218 510048 651454
rect 509728 651134 510048 651218
rect 509728 650898 509770 651134
rect 510006 650898 510048 651134
rect 509728 650866 510048 650898
rect 33568 633454 33888 633486
rect 33568 633218 33610 633454
rect 33846 633218 33888 633454
rect 33568 633134 33888 633218
rect 33568 632898 33610 633134
rect 33846 632898 33888 633134
rect 33568 632866 33888 632898
rect 64288 633454 64608 633486
rect 64288 633218 64330 633454
rect 64566 633218 64608 633454
rect 64288 633134 64608 633218
rect 64288 632898 64330 633134
rect 64566 632898 64608 633134
rect 64288 632866 64608 632898
rect 95008 633454 95328 633486
rect 95008 633218 95050 633454
rect 95286 633218 95328 633454
rect 95008 633134 95328 633218
rect 95008 632898 95050 633134
rect 95286 632898 95328 633134
rect 95008 632866 95328 632898
rect 125728 633454 126048 633486
rect 125728 633218 125770 633454
rect 126006 633218 126048 633454
rect 125728 633134 126048 633218
rect 125728 632898 125770 633134
rect 126006 632898 126048 633134
rect 125728 632866 126048 632898
rect 156448 633454 156768 633486
rect 156448 633218 156490 633454
rect 156726 633218 156768 633454
rect 156448 633134 156768 633218
rect 156448 632898 156490 633134
rect 156726 632898 156768 633134
rect 156448 632866 156768 632898
rect 187168 633454 187488 633486
rect 187168 633218 187210 633454
rect 187446 633218 187488 633454
rect 187168 633134 187488 633218
rect 187168 632898 187210 633134
rect 187446 632898 187488 633134
rect 187168 632866 187488 632898
rect 217888 633454 218208 633486
rect 217888 633218 217930 633454
rect 218166 633218 218208 633454
rect 217888 633134 218208 633218
rect 217888 632898 217930 633134
rect 218166 632898 218208 633134
rect 217888 632866 218208 632898
rect 248608 633454 248928 633486
rect 248608 633218 248650 633454
rect 248886 633218 248928 633454
rect 248608 633134 248928 633218
rect 248608 632898 248650 633134
rect 248886 632898 248928 633134
rect 248608 632866 248928 632898
rect 279328 633454 279648 633486
rect 279328 633218 279370 633454
rect 279606 633218 279648 633454
rect 279328 633134 279648 633218
rect 279328 632898 279370 633134
rect 279606 632898 279648 633134
rect 279328 632866 279648 632898
rect 310048 633454 310368 633486
rect 310048 633218 310090 633454
rect 310326 633218 310368 633454
rect 310048 633134 310368 633218
rect 310048 632898 310090 633134
rect 310326 632898 310368 633134
rect 310048 632866 310368 632898
rect 340768 633454 341088 633486
rect 340768 633218 340810 633454
rect 341046 633218 341088 633454
rect 340768 633134 341088 633218
rect 340768 632898 340810 633134
rect 341046 632898 341088 633134
rect 340768 632866 341088 632898
rect 371488 633454 371808 633486
rect 371488 633218 371530 633454
rect 371766 633218 371808 633454
rect 371488 633134 371808 633218
rect 371488 632898 371530 633134
rect 371766 632898 371808 633134
rect 371488 632866 371808 632898
rect 402208 633454 402528 633486
rect 402208 633218 402250 633454
rect 402486 633218 402528 633454
rect 402208 633134 402528 633218
rect 402208 632898 402250 633134
rect 402486 632898 402528 633134
rect 402208 632866 402528 632898
rect 432928 633454 433248 633486
rect 432928 633218 432970 633454
rect 433206 633218 433248 633454
rect 432928 633134 433248 633218
rect 432928 632898 432970 633134
rect 433206 632898 433248 633134
rect 432928 632866 433248 632898
rect 463648 633454 463968 633486
rect 463648 633218 463690 633454
rect 463926 633218 463968 633454
rect 463648 633134 463968 633218
rect 463648 632898 463690 633134
rect 463926 632898 463968 633134
rect 463648 632866 463968 632898
rect 494368 633454 494688 633486
rect 494368 633218 494410 633454
rect 494646 633218 494688 633454
rect 494368 633134 494688 633218
rect 494368 632898 494410 633134
rect 494646 632898 494688 633134
rect 494368 632866 494688 632898
rect 525088 633454 525408 633486
rect 525088 633218 525130 633454
rect 525366 633218 525408 633454
rect 525088 633134 525408 633218
rect 525088 632898 525130 633134
rect 525366 632898 525408 633134
rect 525088 632866 525408 632898
rect 48928 615454 49248 615486
rect 48928 615218 48970 615454
rect 49206 615218 49248 615454
rect 48928 615134 49248 615218
rect 48928 614898 48970 615134
rect 49206 614898 49248 615134
rect 48928 614866 49248 614898
rect 79648 615454 79968 615486
rect 79648 615218 79690 615454
rect 79926 615218 79968 615454
rect 79648 615134 79968 615218
rect 79648 614898 79690 615134
rect 79926 614898 79968 615134
rect 79648 614866 79968 614898
rect 110368 615454 110688 615486
rect 110368 615218 110410 615454
rect 110646 615218 110688 615454
rect 110368 615134 110688 615218
rect 110368 614898 110410 615134
rect 110646 614898 110688 615134
rect 110368 614866 110688 614898
rect 141088 615454 141408 615486
rect 141088 615218 141130 615454
rect 141366 615218 141408 615454
rect 141088 615134 141408 615218
rect 141088 614898 141130 615134
rect 141366 614898 141408 615134
rect 141088 614866 141408 614898
rect 171808 615454 172128 615486
rect 171808 615218 171850 615454
rect 172086 615218 172128 615454
rect 171808 615134 172128 615218
rect 171808 614898 171850 615134
rect 172086 614898 172128 615134
rect 171808 614866 172128 614898
rect 202528 615454 202848 615486
rect 202528 615218 202570 615454
rect 202806 615218 202848 615454
rect 202528 615134 202848 615218
rect 202528 614898 202570 615134
rect 202806 614898 202848 615134
rect 202528 614866 202848 614898
rect 233248 615454 233568 615486
rect 233248 615218 233290 615454
rect 233526 615218 233568 615454
rect 233248 615134 233568 615218
rect 233248 614898 233290 615134
rect 233526 614898 233568 615134
rect 233248 614866 233568 614898
rect 263968 615454 264288 615486
rect 263968 615218 264010 615454
rect 264246 615218 264288 615454
rect 263968 615134 264288 615218
rect 263968 614898 264010 615134
rect 264246 614898 264288 615134
rect 263968 614866 264288 614898
rect 294688 615454 295008 615486
rect 294688 615218 294730 615454
rect 294966 615218 295008 615454
rect 294688 615134 295008 615218
rect 294688 614898 294730 615134
rect 294966 614898 295008 615134
rect 294688 614866 295008 614898
rect 325408 615454 325728 615486
rect 325408 615218 325450 615454
rect 325686 615218 325728 615454
rect 325408 615134 325728 615218
rect 325408 614898 325450 615134
rect 325686 614898 325728 615134
rect 325408 614866 325728 614898
rect 356128 615454 356448 615486
rect 356128 615218 356170 615454
rect 356406 615218 356448 615454
rect 356128 615134 356448 615218
rect 356128 614898 356170 615134
rect 356406 614898 356448 615134
rect 356128 614866 356448 614898
rect 386848 615454 387168 615486
rect 386848 615218 386890 615454
rect 387126 615218 387168 615454
rect 386848 615134 387168 615218
rect 386848 614898 386890 615134
rect 387126 614898 387168 615134
rect 386848 614866 387168 614898
rect 417568 615454 417888 615486
rect 417568 615218 417610 615454
rect 417846 615218 417888 615454
rect 417568 615134 417888 615218
rect 417568 614898 417610 615134
rect 417846 614898 417888 615134
rect 417568 614866 417888 614898
rect 448288 615454 448608 615486
rect 448288 615218 448330 615454
rect 448566 615218 448608 615454
rect 448288 615134 448608 615218
rect 448288 614898 448330 615134
rect 448566 614898 448608 615134
rect 448288 614866 448608 614898
rect 479008 615454 479328 615486
rect 479008 615218 479050 615454
rect 479286 615218 479328 615454
rect 479008 615134 479328 615218
rect 479008 614898 479050 615134
rect 479286 614898 479328 615134
rect 479008 614866 479328 614898
rect 509728 615454 510048 615486
rect 509728 615218 509770 615454
rect 510006 615218 510048 615454
rect 509728 615134 510048 615218
rect 509728 614898 509770 615134
rect 510006 614898 510048 615134
rect 509728 614866 510048 614898
rect 33568 597454 33888 597486
rect 33568 597218 33610 597454
rect 33846 597218 33888 597454
rect 33568 597134 33888 597218
rect 33568 596898 33610 597134
rect 33846 596898 33888 597134
rect 33568 596866 33888 596898
rect 64288 597454 64608 597486
rect 64288 597218 64330 597454
rect 64566 597218 64608 597454
rect 64288 597134 64608 597218
rect 64288 596898 64330 597134
rect 64566 596898 64608 597134
rect 64288 596866 64608 596898
rect 95008 597454 95328 597486
rect 95008 597218 95050 597454
rect 95286 597218 95328 597454
rect 95008 597134 95328 597218
rect 95008 596898 95050 597134
rect 95286 596898 95328 597134
rect 95008 596866 95328 596898
rect 125728 597454 126048 597486
rect 125728 597218 125770 597454
rect 126006 597218 126048 597454
rect 125728 597134 126048 597218
rect 125728 596898 125770 597134
rect 126006 596898 126048 597134
rect 125728 596866 126048 596898
rect 156448 597454 156768 597486
rect 156448 597218 156490 597454
rect 156726 597218 156768 597454
rect 156448 597134 156768 597218
rect 156448 596898 156490 597134
rect 156726 596898 156768 597134
rect 156448 596866 156768 596898
rect 187168 597454 187488 597486
rect 187168 597218 187210 597454
rect 187446 597218 187488 597454
rect 187168 597134 187488 597218
rect 187168 596898 187210 597134
rect 187446 596898 187488 597134
rect 187168 596866 187488 596898
rect 217888 597454 218208 597486
rect 217888 597218 217930 597454
rect 218166 597218 218208 597454
rect 217888 597134 218208 597218
rect 217888 596898 217930 597134
rect 218166 596898 218208 597134
rect 217888 596866 218208 596898
rect 248608 597454 248928 597486
rect 248608 597218 248650 597454
rect 248886 597218 248928 597454
rect 248608 597134 248928 597218
rect 248608 596898 248650 597134
rect 248886 596898 248928 597134
rect 248608 596866 248928 596898
rect 279328 597454 279648 597486
rect 279328 597218 279370 597454
rect 279606 597218 279648 597454
rect 279328 597134 279648 597218
rect 279328 596898 279370 597134
rect 279606 596898 279648 597134
rect 279328 596866 279648 596898
rect 310048 597454 310368 597486
rect 310048 597218 310090 597454
rect 310326 597218 310368 597454
rect 310048 597134 310368 597218
rect 310048 596898 310090 597134
rect 310326 596898 310368 597134
rect 310048 596866 310368 596898
rect 340768 597454 341088 597486
rect 340768 597218 340810 597454
rect 341046 597218 341088 597454
rect 340768 597134 341088 597218
rect 340768 596898 340810 597134
rect 341046 596898 341088 597134
rect 340768 596866 341088 596898
rect 371488 597454 371808 597486
rect 371488 597218 371530 597454
rect 371766 597218 371808 597454
rect 371488 597134 371808 597218
rect 371488 596898 371530 597134
rect 371766 596898 371808 597134
rect 371488 596866 371808 596898
rect 402208 597454 402528 597486
rect 402208 597218 402250 597454
rect 402486 597218 402528 597454
rect 402208 597134 402528 597218
rect 402208 596898 402250 597134
rect 402486 596898 402528 597134
rect 402208 596866 402528 596898
rect 432928 597454 433248 597486
rect 432928 597218 432970 597454
rect 433206 597218 433248 597454
rect 432928 597134 433248 597218
rect 432928 596898 432970 597134
rect 433206 596898 433248 597134
rect 432928 596866 433248 596898
rect 463648 597454 463968 597486
rect 463648 597218 463690 597454
rect 463926 597218 463968 597454
rect 463648 597134 463968 597218
rect 463648 596898 463690 597134
rect 463926 596898 463968 597134
rect 463648 596866 463968 596898
rect 494368 597454 494688 597486
rect 494368 597218 494410 597454
rect 494646 597218 494688 597454
rect 494368 597134 494688 597218
rect 494368 596898 494410 597134
rect 494646 596898 494688 597134
rect 494368 596866 494688 596898
rect 525088 597454 525408 597486
rect 525088 597218 525130 597454
rect 525366 597218 525408 597454
rect 525088 597134 525408 597218
rect 525088 596898 525130 597134
rect 525366 596898 525408 597134
rect 525088 596866 525408 596898
rect 48928 579454 49248 579486
rect 48928 579218 48970 579454
rect 49206 579218 49248 579454
rect 48928 579134 49248 579218
rect 48928 578898 48970 579134
rect 49206 578898 49248 579134
rect 48928 578866 49248 578898
rect 79648 579454 79968 579486
rect 79648 579218 79690 579454
rect 79926 579218 79968 579454
rect 79648 579134 79968 579218
rect 79648 578898 79690 579134
rect 79926 578898 79968 579134
rect 79648 578866 79968 578898
rect 110368 579454 110688 579486
rect 110368 579218 110410 579454
rect 110646 579218 110688 579454
rect 110368 579134 110688 579218
rect 110368 578898 110410 579134
rect 110646 578898 110688 579134
rect 110368 578866 110688 578898
rect 141088 579454 141408 579486
rect 141088 579218 141130 579454
rect 141366 579218 141408 579454
rect 141088 579134 141408 579218
rect 141088 578898 141130 579134
rect 141366 578898 141408 579134
rect 141088 578866 141408 578898
rect 171808 579454 172128 579486
rect 171808 579218 171850 579454
rect 172086 579218 172128 579454
rect 171808 579134 172128 579218
rect 171808 578898 171850 579134
rect 172086 578898 172128 579134
rect 171808 578866 172128 578898
rect 202528 579454 202848 579486
rect 202528 579218 202570 579454
rect 202806 579218 202848 579454
rect 202528 579134 202848 579218
rect 202528 578898 202570 579134
rect 202806 578898 202848 579134
rect 202528 578866 202848 578898
rect 233248 579454 233568 579486
rect 233248 579218 233290 579454
rect 233526 579218 233568 579454
rect 233248 579134 233568 579218
rect 233248 578898 233290 579134
rect 233526 578898 233568 579134
rect 233248 578866 233568 578898
rect 263968 579454 264288 579486
rect 263968 579218 264010 579454
rect 264246 579218 264288 579454
rect 263968 579134 264288 579218
rect 263968 578898 264010 579134
rect 264246 578898 264288 579134
rect 263968 578866 264288 578898
rect 294688 579454 295008 579486
rect 294688 579218 294730 579454
rect 294966 579218 295008 579454
rect 294688 579134 295008 579218
rect 294688 578898 294730 579134
rect 294966 578898 295008 579134
rect 294688 578866 295008 578898
rect 325408 579454 325728 579486
rect 325408 579218 325450 579454
rect 325686 579218 325728 579454
rect 325408 579134 325728 579218
rect 325408 578898 325450 579134
rect 325686 578898 325728 579134
rect 325408 578866 325728 578898
rect 356128 579454 356448 579486
rect 356128 579218 356170 579454
rect 356406 579218 356448 579454
rect 356128 579134 356448 579218
rect 356128 578898 356170 579134
rect 356406 578898 356448 579134
rect 356128 578866 356448 578898
rect 386848 579454 387168 579486
rect 386848 579218 386890 579454
rect 387126 579218 387168 579454
rect 386848 579134 387168 579218
rect 386848 578898 386890 579134
rect 387126 578898 387168 579134
rect 386848 578866 387168 578898
rect 417568 579454 417888 579486
rect 417568 579218 417610 579454
rect 417846 579218 417888 579454
rect 417568 579134 417888 579218
rect 417568 578898 417610 579134
rect 417846 578898 417888 579134
rect 417568 578866 417888 578898
rect 448288 579454 448608 579486
rect 448288 579218 448330 579454
rect 448566 579218 448608 579454
rect 448288 579134 448608 579218
rect 448288 578898 448330 579134
rect 448566 578898 448608 579134
rect 448288 578866 448608 578898
rect 479008 579454 479328 579486
rect 479008 579218 479050 579454
rect 479286 579218 479328 579454
rect 479008 579134 479328 579218
rect 479008 578898 479050 579134
rect 479286 578898 479328 579134
rect 479008 578866 479328 578898
rect 509728 579454 510048 579486
rect 509728 579218 509770 579454
rect 510006 579218 510048 579454
rect 509728 579134 510048 579218
rect 509728 578898 509770 579134
rect 510006 578898 510048 579134
rect 509728 578866 510048 578898
rect 33568 561454 33888 561486
rect 33568 561218 33610 561454
rect 33846 561218 33888 561454
rect 33568 561134 33888 561218
rect 33568 560898 33610 561134
rect 33846 560898 33888 561134
rect 33568 560866 33888 560898
rect 64288 561454 64608 561486
rect 64288 561218 64330 561454
rect 64566 561218 64608 561454
rect 64288 561134 64608 561218
rect 64288 560898 64330 561134
rect 64566 560898 64608 561134
rect 64288 560866 64608 560898
rect 95008 561454 95328 561486
rect 95008 561218 95050 561454
rect 95286 561218 95328 561454
rect 95008 561134 95328 561218
rect 95008 560898 95050 561134
rect 95286 560898 95328 561134
rect 95008 560866 95328 560898
rect 125728 561454 126048 561486
rect 125728 561218 125770 561454
rect 126006 561218 126048 561454
rect 125728 561134 126048 561218
rect 125728 560898 125770 561134
rect 126006 560898 126048 561134
rect 125728 560866 126048 560898
rect 156448 561454 156768 561486
rect 156448 561218 156490 561454
rect 156726 561218 156768 561454
rect 156448 561134 156768 561218
rect 156448 560898 156490 561134
rect 156726 560898 156768 561134
rect 156448 560866 156768 560898
rect 187168 561454 187488 561486
rect 187168 561218 187210 561454
rect 187446 561218 187488 561454
rect 187168 561134 187488 561218
rect 187168 560898 187210 561134
rect 187446 560898 187488 561134
rect 187168 560866 187488 560898
rect 217888 561454 218208 561486
rect 217888 561218 217930 561454
rect 218166 561218 218208 561454
rect 217888 561134 218208 561218
rect 217888 560898 217930 561134
rect 218166 560898 218208 561134
rect 217888 560866 218208 560898
rect 248608 561454 248928 561486
rect 248608 561218 248650 561454
rect 248886 561218 248928 561454
rect 248608 561134 248928 561218
rect 248608 560898 248650 561134
rect 248886 560898 248928 561134
rect 248608 560866 248928 560898
rect 279328 561454 279648 561486
rect 279328 561218 279370 561454
rect 279606 561218 279648 561454
rect 279328 561134 279648 561218
rect 279328 560898 279370 561134
rect 279606 560898 279648 561134
rect 279328 560866 279648 560898
rect 310048 561454 310368 561486
rect 310048 561218 310090 561454
rect 310326 561218 310368 561454
rect 310048 561134 310368 561218
rect 310048 560898 310090 561134
rect 310326 560898 310368 561134
rect 310048 560866 310368 560898
rect 340768 561454 341088 561486
rect 340768 561218 340810 561454
rect 341046 561218 341088 561454
rect 340768 561134 341088 561218
rect 340768 560898 340810 561134
rect 341046 560898 341088 561134
rect 340768 560866 341088 560898
rect 371488 561454 371808 561486
rect 371488 561218 371530 561454
rect 371766 561218 371808 561454
rect 371488 561134 371808 561218
rect 371488 560898 371530 561134
rect 371766 560898 371808 561134
rect 371488 560866 371808 560898
rect 402208 561454 402528 561486
rect 402208 561218 402250 561454
rect 402486 561218 402528 561454
rect 402208 561134 402528 561218
rect 402208 560898 402250 561134
rect 402486 560898 402528 561134
rect 402208 560866 402528 560898
rect 432928 561454 433248 561486
rect 432928 561218 432970 561454
rect 433206 561218 433248 561454
rect 432928 561134 433248 561218
rect 432928 560898 432970 561134
rect 433206 560898 433248 561134
rect 432928 560866 433248 560898
rect 463648 561454 463968 561486
rect 463648 561218 463690 561454
rect 463926 561218 463968 561454
rect 463648 561134 463968 561218
rect 463648 560898 463690 561134
rect 463926 560898 463968 561134
rect 463648 560866 463968 560898
rect 494368 561454 494688 561486
rect 494368 561218 494410 561454
rect 494646 561218 494688 561454
rect 494368 561134 494688 561218
rect 494368 560898 494410 561134
rect 494646 560898 494688 561134
rect 494368 560866 494688 560898
rect 525088 561454 525408 561486
rect 525088 561218 525130 561454
rect 525366 561218 525408 561454
rect 525088 561134 525408 561218
rect 525088 560898 525130 561134
rect 525366 560898 525408 561134
rect 525088 560866 525408 560898
rect 48928 543454 49248 543486
rect 48928 543218 48970 543454
rect 49206 543218 49248 543454
rect 48928 543134 49248 543218
rect 48928 542898 48970 543134
rect 49206 542898 49248 543134
rect 48928 542866 49248 542898
rect 79648 543454 79968 543486
rect 79648 543218 79690 543454
rect 79926 543218 79968 543454
rect 79648 543134 79968 543218
rect 79648 542898 79690 543134
rect 79926 542898 79968 543134
rect 79648 542866 79968 542898
rect 110368 543454 110688 543486
rect 110368 543218 110410 543454
rect 110646 543218 110688 543454
rect 110368 543134 110688 543218
rect 110368 542898 110410 543134
rect 110646 542898 110688 543134
rect 110368 542866 110688 542898
rect 141088 543454 141408 543486
rect 141088 543218 141130 543454
rect 141366 543218 141408 543454
rect 141088 543134 141408 543218
rect 141088 542898 141130 543134
rect 141366 542898 141408 543134
rect 141088 542866 141408 542898
rect 171808 543454 172128 543486
rect 171808 543218 171850 543454
rect 172086 543218 172128 543454
rect 171808 543134 172128 543218
rect 171808 542898 171850 543134
rect 172086 542898 172128 543134
rect 171808 542866 172128 542898
rect 202528 543454 202848 543486
rect 202528 543218 202570 543454
rect 202806 543218 202848 543454
rect 202528 543134 202848 543218
rect 202528 542898 202570 543134
rect 202806 542898 202848 543134
rect 202528 542866 202848 542898
rect 233248 543454 233568 543486
rect 233248 543218 233290 543454
rect 233526 543218 233568 543454
rect 233248 543134 233568 543218
rect 233248 542898 233290 543134
rect 233526 542898 233568 543134
rect 233248 542866 233568 542898
rect 263968 543454 264288 543486
rect 263968 543218 264010 543454
rect 264246 543218 264288 543454
rect 263968 543134 264288 543218
rect 263968 542898 264010 543134
rect 264246 542898 264288 543134
rect 263968 542866 264288 542898
rect 294688 543454 295008 543486
rect 294688 543218 294730 543454
rect 294966 543218 295008 543454
rect 294688 543134 295008 543218
rect 294688 542898 294730 543134
rect 294966 542898 295008 543134
rect 294688 542866 295008 542898
rect 325408 543454 325728 543486
rect 325408 543218 325450 543454
rect 325686 543218 325728 543454
rect 325408 543134 325728 543218
rect 325408 542898 325450 543134
rect 325686 542898 325728 543134
rect 325408 542866 325728 542898
rect 356128 543454 356448 543486
rect 356128 543218 356170 543454
rect 356406 543218 356448 543454
rect 356128 543134 356448 543218
rect 356128 542898 356170 543134
rect 356406 542898 356448 543134
rect 356128 542866 356448 542898
rect 386848 543454 387168 543486
rect 386848 543218 386890 543454
rect 387126 543218 387168 543454
rect 386848 543134 387168 543218
rect 386848 542898 386890 543134
rect 387126 542898 387168 543134
rect 386848 542866 387168 542898
rect 417568 543454 417888 543486
rect 417568 543218 417610 543454
rect 417846 543218 417888 543454
rect 417568 543134 417888 543218
rect 417568 542898 417610 543134
rect 417846 542898 417888 543134
rect 417568 542866 417888 542898
rect 448288 543454 448608 543486
rect 448288 543218 448330 543454
rect 448566 543218 448608 543454
rect 448288 543134 448608 543218
rect 448288 542898 448330 543134
rect 448566 542898 448608 543134
rect 448288 542866 448608 542898
rect 479008 543454 479328 543486
rect 479008 543218 479050 543454
rect 479286 543218 479328 543454
rect 479008 543134 479328 543218
rect 479008 542898 479050 543134
rect 479286 542898 479328 543134
rect 479008 542866 479328 542898
rect 509728 543454 510048 543486
rect 509728 543218 509770 543454
rect 510006 543218 510048 543454
rect 509728 543134 510048 543218
rect 509728 542898 509770 543134
rect 510006 542898 510048 543134
rect 509728 542866 510048 542898
rect 33568 525454 33888 525486
rect 33568 525218 33610 525454
rect 33846 525218 33888 525454
rect 33568 525134 33888 525218
rect 33568 524898 33610 525134
rect 33846 524898 33888 525134
rect 33568 524866 33888 524898
rect 64288 525454 64608 525486
rect 64288 525218 64330 525454
rect 64566 525218 64608 525454
rect 64288 525134 64608 525218
rect 64288 524898 64330 525134
rect 64566 524898 64608 525134
rect 64288 524866 64608 524898
rect 95008 525454 95328 525486
rect 95008 525218 95050 525454
rect 95286 525218 95328 525454
rect 95008 525134 95328 525218
rect 95008 524898 95050 525134
rect 95286 524898 95328 525134
rect 95008 524866 95328 524898
rect 125728 525454 126048 525486
rect 125728 525218 125770 525454
rect 126006 525218 126048 525454
rect 125728 525134 126048 525218
rect 125728 524898 125770 525134
rect 126006 524898 126048 525134
rect 125728 524866 126048 524898
rect 156448 525454 156768 525486
rect 156448 525218 156490 525454
rect 156726 525218 156768 525454
rect 156448 525134 156768 525218
rect 156448 524898 156490 525134
rect 156726 524898 156768 525134
rect 156448 524866 156768 524898
rect 187168 525454 187488 525486
rect 187168 525218 187210 525454
rect 187446 525218 187488 525454
rect 187168 525134 187488 525218
rect 187168 524898 187210 525134
rect 187446 524898 187488 525134
rect 187168 524866 187488 524898
rect 217888 525454 218208 525486
rect 217888 525218 217930 525454
rect 218166 525218 218208 525454
rect 217888 525134 218208 525218
rect 217888 524898 217930 525134
rect 218166 524898 218208 525134
rect 217888 524866 218208 524898
rect 248608 525454 248928 525486
rect 248608 525218 248650 525454
rect 248886 525218 248928 525454
rect 248608 525134 248928 525218
rect 248608 524898 248650 525134
rect 248886 524898 248928 525134
rect 248608 524866 248928 524898
rect 279328 525454 279648 525486
rect 279328 525218 279370 525454
rect 279606 525218 279648 525454
rect 279328 525134 279648 525218
rect 279328 524898 279370 525134
rect 279606 524898 279648 525134
rect 279328 524866 279648 524898
rect 310048 525454 310368 525486
rect 310048 525218 310090 525454
rect 310326 525218 310368 525454
rect 310048 525134 310368 525218
rect 310048 524898 310090 525134
rect 310326 524898 310368 525134
rect 310048 524866 310368 524898
rect 340768 525454 341088 525486
rect 340768 525218 340810 525454
rect 341046 525218 341088 525454
rect 340768 525134 341088 525218
rect 340768 524898 340810 525134
rect 341046 524898 341088 525134
rect 340768 524866 341088 524898
rect 371488 525454 371808 525486
rect 371488 525218 371530 525454
rect 371766 525218 371808 525454
rect 371488 525134 371808 525218
rect 371488 524898 371530 525134
rect 371766 524898 371808 525134
rect 371488 524866 371808 524898
rect 402208 525454 402528 525486
rect 402208 525218 402250 525454
rect 402486 525218 402528 525454
rect 402208 525134 402528 525218
rect 402208 524898 402250 525134
rect 402486 524898 402528 525134
rect 402208 524866 402528 524898
rect 432928 525454 433248 525486
rect 432928 525218 432970 525454
rect 433206 525218 433248 525454
rect 432928 525134 433248 525218
rect 432928 524898 432970 525134
rect 433206 524898 433248 525134
rect 432928 524866 433248 524898
rect 463648 525454 463968 525486
rect 463648 525218 463690 525454
rect 463926 525218 463968 525454
rect 463648 525134 463968 525218
rect 463648 524898 463690 525134
rect 463926 524898 463968 525134
rect 463648 524866 463968 524898
rect 494368 525454 494688 525486
rect 494368 525218 494410 525454
rect 494646 525218 494688 525454
rect 494368 525134 494688 525218
rect 494368 524898 494410 525134
rect 494646 524898 494688 525134
rect 494368 524866 494688 524898
rect 525088 525454 525408 525486
rect 525088 525218 525130 525454
rect 525366 525218 525408 525454
rect 525088 525134 525408 525218
rect 525088 524898 525130 525134
rect 525366 524898 525408 525134
rect 525088 524866 525408 524898
rect 48928 507454 49248 507486
rect 48928 507218 48970 507454
rect 49206 507218 49248 507454
rect 48928 507134 49248 507218
rect 48928 506898 48970 507134
rect 49206 506898 49248 507134
rect 48928 506866 49248 506898
rect 79648 507454 79968 507486
rect 79648 507218 79690 507454
rect 79926 507218 79968 507454
rect 79648 507134 79968 507218
rect 79648 506898 79690 507134
rect 79926 506898 79968 507134
rect 79648 506866 79968 506898
rect 110368 507454 110688 507486
rect 110368 507218 110410 507454
rect 110646 507218 110688 507454
rect 110368 507134 110688 507218
rect 110368 506898 110410 507134
rect 110646 506898 110688 507134
rect 110368 506866 110688 506898
rect 141088 507454 141408 507486
rect 141088 507218 141130 507454
rect 141366 507218 141408 507454
rect 141088 507134 141408 507218
rect 141088 506898 141130 507134
rect 141366 506898 141408 507134
rect 141088 506866 141408 506898
rect 171808 507454 172128 507486
rect 171808 507218 171850 507454
rect 172086 507218 172128 507454
rect 171808 507134 172128 507218
rect 171808 506898 171850 507134
rect 172086 506898 172128 507134
rect 171808 506866 172128 506898
rect 202528 507454 202848 507486
rect 202528 507218 202570 507454
rect 202806 507218 202848 507454
rect 202528 507134 202848 507218
rect 202528 506898 202570 507134
rect 202806 506898 202848 507134
rect 202528 506866 202848 506898
rect 233248 507454 233568 507486
rect 233248 507218 233290 507454
rect 233526 507218 233568 507454
rect 233248 507134 233568 507218
rect 233248 506898 233290 507134
rect 233526 506898 233568 507134
rect 233248 506866 233568 506898
rect 263968 507454 264288 507486
rect 263968 507218 264010 507454
rect 264246 507218 264288 507454
rect 263968 507134 264288 507218
rect 263968 506898 264010 507134
rect 264246 506898 264288 507134
rect 263968 506866 264288 506898
rect 294688 507454 295008 507486
rect 294688 507218 294730 507454
rect 294966 507218 295008 507454
rect 294688 507134 295008 507218
rect 294688 506898 294730 507134
rect 294966 506898 295008 507134
rect 294688 506866 295008 506898
rect 325408 507454 325728 507486
rect 325408 507218 325450 507454
rect 325686 507218 325728 507454
rect 325408 507134 325728 507218
rect 325408 506898 325450 507134
rect 325686 506898 325728 507134
rect 325408 506866 325728 506898
rect 356128 507454 356448 507486
rect 356128 507218 356170 507454
rect 356406 507218 356448 507454
rect 356128 507134 356448 507218
rect 356128 506898 356170 507134
rect 356406 506898 356448 507134
rect 356128 506866 356448 506898
rect 386848 507454 387168 507486
rect 386848 507218 386890 507454
rect 387126 507218 387168 507454
rect 386848 507134 387168 507218
rect 386848 506898 386890 507134
rect 387126 506898 387168 507134
rect 386848 506866 387168 506898
rect 417568 507454 417888 507486
rect 417568 507218 417610 507454
rect 417846 507218 417888 507454
rect 417568 507134 417888 507218
rect 417568 506898 417610 507134
rect 417846 506898 417888 507134
rect 417568 506866 417888 506898
rect 448288 507454 448608 507486
rect 448288 507218 448330 507454
rect 448566 507218 448608 507454
rect 448288 507134 448608 507218
rect 448288 506898 448330 507134
rect 448566 506898 448608 507134
rect 448288 506866 448608 506898
rect 479008 507454 479328 507486
rect 479008 507218 479050 507454
rect 479286 507218 479328 507454
rect 479008 507134 479328 507218
rect 479008 506898 479050 507134
rect 479286 506898 479328 507134
rect 479008 506866 479328 506898
rect 509728 507454 510048 507486
rect 509728 507218 509770 507454
rect 510006 507218 510048 507454
rect 509728 507134 510048 507218
rect 509728 506898 509770 507134
rect 510006 506898 510048 507134
rect 509728 506866 510048 506898
rect 33568 489454 33888 489486
rect 33568 489218 33610 489454
rect 33846 489218 33888 489454
rect 33568 489134 33888 489218
rect 33568 488898 33610 489134
rect 33846 488898 33888 489134
rect 33568 488866 33888 488898
rect 64288 489454 64608 489486
rect 64288 489218 64330 489454
rect 64566 489218 64608 489454
rect 64288 489134 64608 489218
rect 64288 488898 64330 489134
rect 64566 488898 64608 489134
rect 64288 488866 64608 488898
rect 95008 489454 95328 489486
rect 95008 489218 95050 489454
rect 95286 489218 95328 489454
rect 95008 489134 95328 489218
rect 95008 488898 95050 489134
rect 95286 488898 95328 489134
rect 95008 488866 95328 488898
rect 125728 489454 126048 489486
rect 125728 489218 125770 489454
rect 126006 489218 126048 489454
rect 125728 489134 126048 489218
rect 125728 488898 125770 489134
rect 126006 488898 126048 489134
rect 125728 488866 126048 488898
rect 156448 489454 156768 489486
rect 156448 489218 156490 489454
rect 156726 489218 156768 489454
rect 156448 489134 156768 489218
rect 156448 488898 156490 489134
rect 156726 488898 156768 489134
rect 156448 488866 156768 488898
rect 187168 489454 187488 489486
rect 187168 489218 187210 489454
rect 187446 489218 187488 489454
rect 187168 489134 187488 489218
rect 187168 488898 187210 489134
rect 187446 488898 187488 489134
rect 187168 488866 187488 488898
rect 217888 489454 218208 489486
rect 217888 489218 217930 489454
rect 218166 489218 218208 489454
rect 217888 489134 218208 489218
rect 217888 488898 217930 489134
rect 218166 488898 218208 489134
rect 217888 488866 218208 488898
rect 248608 489454 248928 489486
rect 248608 489218 248650 489454
rect 248886 489218 248928 489454
rect 248608 489134 248928 489218
rect 248608 488898 248650 489134
rect 248886 488898 248928 489134
rect 248608 488866 248928 488898
rect 279328 489454 279648 489486
rect 279328 489218 279370 489454
rect 279606 489218 279648 489454
rect 279328 489134 279648 489218
rect 279328 488898 279370 489134
rect 279606 488898 279648 489134
rect 279328 488866 279648 488898
rect 310048 489454 310368 489486
rect 310048 489218 310090 489454
rect 310326 489218 310368 489454
rect 310048 489134 310368 489218
rect 310048 488898 310090 489134
rect 310326 488898 310368 489134
rect 310048 488866 310368 488898
rect 340768 489454 341088 489486
rect 340768 489218 340810 489454
rect 341046 489218 341088 489454
rect 340768 489134 341088 489218
rect 340768 488898 340810 489134
rect 341046 488898 341088 489134
rect 340768 488866 341088 488898
rect 371488 489454 371808 489486
rect 371488 489218 371530 489454
rect 371766 489218 371808 489454
rect 371488 489134 371808 489218
rect 371488 488898 371530 489134
rect 371766 488898 371808 489134
rect 371488 488866 371808 488898
rect 402208 489454 402528 489486
rect 402208 489218 402250 489454
rect 402486 489218 402528 489454
rect 402208 489134 402528 489218
rect 402208 488898 402250 489134
rect 402486 488898 402528 489134
rect 402208 488866 402528 488898
rect 432928 489454 433248 489486
rect 432928 489218 432970 489454
rect 433206 489218 433248 489454
rect 432928 489134 433248 489218
rect 432928 488898 432970 489134
rect 433206 488898 433248 489134
rect 432928 488866 433248 488898
rect 463648 489454 463968 489486
rect 463648 489218 463690 489454
rect 463926 489218 463968 489454
rect 463648 489134 463968 489218
rect 463648 488898 463690 489134
rect 463926 488898 463968 489134
rect 463648 488866 463968 488898
rect 494368 489454 494688 489486
rect 494368 489218 494410 489454
rect 494646 489218 494688 489454
rect 494368 489134 494688 489218
rect 494368 488898 494410 489134
rect 494646 488898 494688 489134
rect 494368 488866 494688 488898
rect 525088 489454 525408 489486
rect 525088 489218 525130 489454
rect 525366 489218 525408 489454
rect 525088 489134 525408 489218
rect 525088 488898 525130 489134
rect 525366 488898 525408 489134
rect 525088 488866 525408 488898
rect 48928 471454 49248 471486
rect 48928 471218 48970 471454
rect 49206 471218 49248 471454
rect 48928 471134 49248 471218
rect 48928 470898 48970 471134
rect 49206 470898 49248 471134
rect 48928 470866 49248 470898
rect 79648 471454 79968 471486
rect 79648 471218 79690 471454
rect 79926 471218 79968 471454
rect 79648 471134 79968 471218
rect 79648 470898 79690 471134
rect 79926 470898 79968 471134
rect 79648 470866 79968 470898
rect 110368 471454 110688 471486
rect 110368 471218 110410 471454
rect 110646 471218 110688 471454
rect 110368 471134 110688 471218
rect 110368 470898 110410 471134
rect 110646 470898 110688 471134
rect 110368 470866 110688 470898
rect 141088 471454 141408 471486
rect 141088 471218 141130 471454
rect 141366 471218 141408 471454
rect 141088 471134 141408 471218
rect 141088 470898 141130 471134
rect 141366 470898 141408 471134
rect 141088 470866 141408 470898
rect 171808 471454 172128 471486
rect 171808 471218 171850 471454
rect 172086 471218 172128 471454
rect 171808 471134 172128 471218
rect 171808 470898 171850 471134
rect 172086 470898 172128 471134
rect 171808 470866 172128 470898
rect 202528 471454 202848 471486
rect 202528 471218 202570 471454
rect 202806 471218 202848 471454
rect 202528 471134 202848 471218
rect 202528 470898 202570 471134
rect 202806 470898 202848 471134
rect 202528 470866 202848 470898
rect 233248 471454 233568 471486
rect 233248 471218 233290 471454
rect 233526 471218 233568 471454
rect 233248 471134 233568 471218
rect 233248 470898 233290 471134
rect 233526 470898 233568 471134
rect 233248 470866 233568 470898
rect 263968 471454 264288 471486
rect 263968 471218 264010 471454
rect 264246 471218 264288 471454
rect 263968 471134 264288 471218
rect 263968 470898 264010 471134
rect 264246 470898 264288 471134
rect 263968 470866 264288 470898
rect 294688 471454 295008 471486
rect 294688 471218 294730 471454
rect 294966 471218 295008 471454
rect 294688 471134 295008 471218
rect 294688 470898 294730 471134
rect 294966 470898 295008 471134
rect 294688 470866 295008 470898
rect 325408 471454 325728 471486
rect 325408 471218 325450 471454
rect 325686 471218 325728 471454
rect 325408 471134 325728 471218
rect 325408 470898 325450 471134
rect 325686 470898 325728 471134
rect 325408 470866 325728 470898
rect 356128 471454 356448 471486
rect 356128 471218 356170 471454
rect 356406 471218 356448 471454
rect 356128 471134 356448 471218
rect 356128 470898 356170 471134
rect 356406 470898 356448 471134
rect 356128 470866 356448 470898
rect 386848 471454 387168 471486
rect 386848 471218 386890 471454
rect 387126 471218 387168 471454
rect 386848 471134 387168 471218
rect 386848 470898 386890 471134
rect 387126 470898 387168 471134
rect 386848 470866 387168 470898
rect 417568 471454 417888 471486
rect 417568 471218 417610 471454
rect 417846 471218 417888 471454
rect 417568 471134 417888 471218
rect 417568 470898 417610 471134
rect 417846 470898 417888 471134
rect 417568 470866 417888 470898
rect 448288 471454 448608 471486
rect 448288 471218 448330 471454
rect 448566 471218 448608 471454
rect 448288 471134 448608 471218
rect 448288 470898 448330 471134
rect 448566 470898 448608 471134
rect 448288 470866 448608 470898
rect 479008 471454 479328 471486
rect 479008 471218 479050 471454
rect 479286 471218 479328 471454
rect 479008 471134 479328 471218
rect 479008 470898 479050 471134
rect 479286 470898 479328 471134
rect 479008 470866 479328 470898
rect 509728 471454 510048 471486
rect 509728 471218 509770 471454
rect 510006 471218 510048 471454
rect 509728 471134 510048 471218
rect 509728 470898 509770 471134
rect 510006 470898 510048 471134
rect 509728 470866 510048 470898
rect 33568 453454 33888 453486
rect 33568 453218 33610 453454
rect 33846 453218 33888 453454
rect 33568 453134 33888 453218
rect 33568 452898 33610 453134
rect 33846 452898 33888 453134
rect 33568 452866 33888 452898
rect 64288 453454 64608 453486
rect 64288 453218 64330 453454
rect 64566 453218 64608 453454
rect 64288 453134 64608 453218
rect 64288 452898 64330 453134
rect 64566 452898 64608 453134
rect 64288 452866 64608 452898
rect 95008 453454 95328 453486
rect 95008 453218 95050 453454
rect 95286 453218 95328 453454
rect 95008 453134 95328 453218
rect 95008 452898 95050 453134
rect 95286 452898 95328 453134
rect 95008 452866 95328 452898
rect 125728 453454 126048 453486
rect 125728 453218 125770 453454
rect 126006 453218 126048 453454
rect 125728 453134 126048 453218
rect 125728 452898 125770 453134
rect 126006 452898 126048 453134
rect 125728 452866 126048 452898
rect 156448 453454 156768 453486
rect 156448 453218 156490 453454
rect 156726 453218 156768 453454
rect 156448 453134 156768 453218
rect 156448 452898 156490 453134
rect 156726 452898 156768 453134
rect 156448 452866 156768 452898
rect 187168 453454 187488 453486
rect 187168 453218 187210 453454
rect 187446 453218 187488 453454
rect 187168 453134 187488 453218
rect 187168 452898 187210 453134
rect 187446 452898 187488 453134
rect 187168 452866 187488 452898
rect 217888 453454 218208 453486
rect 217888 453218 217930 453454
rect 218166 453218 218208 453454
rect 217888 453134 218208 453218
rect 217888 452898 217930 453134
rect 218166 452898 218208 453134
rect 217888 452866 218208 452898
rect 248608 453454 248928 453486
rect 248608 453218 248650 453454
rect 248886 453218 248928 453454
rect 248608 453134 248928 453218
rect 248608 452898 248650 453134
rect 248886 452898 248928 453134
rect 248608 452866 248928 452898
rect 279328 453454 279648 453486
rect 279328 453218 279370 453454
rect 279606 453218 279648 453454
rect 279328 453134 279648 453218
rect 279328 452898 279370 453134
rect 279606 452898 279648 453134
rect 279328 452866 279648 452898
rect 310048 453454 310368 453486
rect 310048 453218 310090 453454
rect 310326 453218 310368 453454
rect 310048 453134 310368 453218
rect 310048 452898 310090 453134
rect 310326 452898 310368 453134
rect 310048 452866 310368 452898
rect 340768 453454 341088 453486
rect 340768 453218 340810 453454
rect 341046 453218 341088 453454
rect 340768 453134 341088 453218
rect 340768 452898 340810 453134
rect 341046 452898 341088 453134
rect 340768 452866 341088 452898
rect 371488 453454 371808 453486
rect 371488 453218 371530 453454
rect 371766 453218 371808 453454
rect 371488 453134 371808 453218
rect 371488 452898 371530 453134
rect 371766 452898 371808 453134
rect 371488 452866 371808 452898
rect 402208 453454 402528 453486
rect 402208 453218 402250 453454
rect 402486 453218 402528 453454
rect 402208 453134 402528 453218
rect 402208 452898 402250 453134
rect 402486 452898 402528 453134
rect 402208 452866 402528 452898
rect 432928 453454 433248 453486
rect 432928 453218 432970 453454
rect 433206 453218 433248 453454
rect 432928 453134 433248 453218
rect 432928 452898 432970 453134
rect 433206 452898 433248 453134
rect 432928 452866 433248 452898
rect 463648 453454 463968 453486
rect 463648 453218 463690 453454
rect 463926 453218 463968 453454
rect 463648 453134 463968 453218
rect 463648 452898 463690 453134
rect 463926 452898 463968 453134
rect 463648 452866 463968 452898
rect 494368 453454 494688 453486
rect 494368 453218 494410 453454
rect 494646 453218 494688 453454
rect 494368 453134 494688 453218
rect 494368 452898 494410 453134
rect 494646 452898 494688 453134
rect 494368 452866 494688 452898
rect 525088 453454 525408 453486
rect 525088 453218 525130 453454
rect 525366 453218 525408 453454
rect 525088 453134 525408 453218
rect 525088 452898 525130 453134
rect 525366 452898 525408 453134
rect 525088 452866 525408 452898
rect 48928 435454 49248 435486
rect 48928 435218 48970 435454
rect 49206 435218 49248 435454
rect 48928 435134 49248 435218
rect 48928 434898 48970 435134
rect 49206 434898 49248 435134
rect 48928 434866 49248 434898
rect 79648 435454 79968 435486
rect 79648 435218 79690 435454
rect 79926 435218 79968 435454
rect 79648 435134 79968 435218
rect 79648 434898 79690 435134
rect 79926 434898 79968 435134
rect 79648 434866 79968 434898
rect 110368 435454 110688 435486
rect 110368 435218 110410 435454
rect 110646 435218 110688 435454
rect 110368 435134 110688 435218
rect 110368 434898 110410 435134
rect 110646 434898 110688 435134
rect 110368 434866 110688 434898
rect 141088 435454 141408 435486
rect 141088 435218 141130 435454
rect 141366 435218 141408 435454
rect 141088 435134 141408 435218
rect 141088 434898 141130 435134
rect 141366 434898 141408 435134
rect 141088 434866 141408 434898
rect 171808 435454 172128 435486
rect 171808 435218 171850 435454
rect 172086 435218 172128 435454
rect 171808 435134 172128 435218
rect 171808 434898 171850 435134
rect 172086 434898 172128 435134
rect 171808 434866 172128 434898
rect 202528 435454 202848 435486
rect 202528 435218 202570 435454
rect 202806 435218 202848 435454
rect 202528 435134 202848 435218
rect 202528 434898 202570 435134
rect 202806 434898 202848 435134
rect 202528 434866 202848 434898
rect 233248 435454 233568 435486
rect 233248 435218 233290 435454
rect 233526 435218 233568 435454
rect 233248 435134 233568 435218
rect 233248 434898 233290 435134
rect 233526 434898 233568 435134
rect 233248 434866 233568 434898
rect 263968 435454 264288 435486
rect 263968 435218 264010 435454
rect 264246 435218 264288 435454
rect 263968 435134 264288 435218
rect 263968 434898 264010 435134
rect 264246 434898 264288 435134
rect 263968 434866 264288 434898
rect 294688 435454 295008 435486
rect 294688 435218 294730 435454
rect 294966 435218 295008 435454
rect 294688 435134 295008 435218
rect 294688 434898 294730 435134
rect 294966 434898 295008 435134
rect 294688 434866 295008 434898
rect 325408 435454 325728 435486
rect 325408 435218 325450 435454
rect 325686 435218 325728 435454
rect 325408 435134 325728 435218
rect 325408 434898 325450 435134
rect 325686 434898 325728 435134
rect 325408 434866 325728 434898
rect 356128 435454 356448 435486
rect 356128 435218 356170 435454
rect 356406 435218 356448 435454
rect 356128 435134 356448 435218
rect 356128 434898 356170 435134
rect 356406 434898 356448 435134
rect 356128 434866 356448 434898
rect 386848 435454 387168 435486
rect 386848 435218 386890 435454
rect 387126 435218 387168 435454
rect 386848 435134 387168 435218
rect 386848 434898 386890 435134
rect 387126 434898 387168 435134
rect 386848 434866 387168 434898
rect 417568 435454 417888 435486
rect 417568 435218 417610 435454
rect 417846 435218 417888 435454
rect 417568 435134 417888 435218
rect 417568 434898 417610 435134
rect 417846 434898 417888 435134
rect 417568 434866 417888 434898
rect 448288 435454 448608 435486
rect 448288 435218 448330 435454
rect 448566 435218 448608 435454
rect 448288 435134 448608 435218
rect 448288 434898 448330 435134
rect 448566 434898 448608 435134
rect 448288 434866 448608 434898
rect 479008 435454 479328 435486
rect 479008 435218 479050 435454
rect 479286 435218 479328 435454
rect 479008 435134 479328 435218
rect 479008 434898 479050 435134
rect 479286 434898 479328 435134
rect 479008 434866 479328 434898
rect 509728 435454 510048 435486
rect 509728 435218 509770 435454
rect 510006 435218 510048 435454
rect 509728 435134 510048 435218
rect 509728 434898 509770 435134
rect 510006 434898 510048 435134
rect 509728 434866 510048 434898
rect 33568 417454 33888 417486
rect 33568 417218 33610 417454
rect 33846 417218 33888 417454
rect 33568 417134 33888 417218
rect 33568 416898 33610 417134
rect 33846 416898 33888 417134
rect 33568 416866 33888 416898
rect 64288 417454 64608 417486
rect 64288 417218 64330 417454
rect 64566 417218 64608 417454
rect 64288 417134 64608 417218
rect 64288 416898 64330 417134
rect 64566 416898 64608 417134
rect 64288 416866 64608 416898
rect 95008 417454 95328 417486
rect 95008 417218 95050 417454
rect 95286 417218 95328 417454
rect 95008 417134 95328 417218
rect 95008 416898 95050 417134
rect 95286 416898 95328 417134
rect 95008 416866 95328 416898
rect 125728 417454 126048 417486
rect 125728 417218 125770 417454
rect 126006 417218 126048 417454
rect 125728 417134 126048 417218
rect 125728 416898 125770 417134
rect 126006 416898 126048 417134
rect 125728 416866 126048 416898
rect 156448 417454 156768 417486
rect 156448 417218 156490 417454
rect 156726 417218 156768 417454
rect 156448 417134 156768 417218
rect 156448 416898 156490 417134
rect 156726 416898 156768 417134
rect 156448 416866 156768 416898
rect 187168 417454 187488 417486
rect 187168 417218 187210 417454
rect 187446 417218 187488 417454
rect 187168 417134 187488 417218
rect 187168 416898 187210 417134
rect 187446 416898 187488 417134
rect 187168 416866 187488 416898
rect 217888 417454 218208 417486
rect 217888 417218 217930 417454
rect 218166 417218 218208 417454
rect 217888 417134 218208 417218
rect 217888 416898 217930 417134
rect 218166 416898 218208 417134
rect 217888 416866 218208 416898
rect 248608 417454 248928 417486
rect 248608 417218 248650 417454
rect 248886 417218 248928 417454
rect 248608 417134 248928 417218
rect 248608 416898 248650 417134
rect 248886 416898 248928 417134
rect 248608 416866 248928 416898
rect 279328 417454 279648 417486
rect 279328 417218 279370 417454
rect 279606 417218 279648 417454
rect 279328 417134 279648 417218
rect 279328 416898 279370 417134
rect 279606 416898 279648 417134
rect 279328 416866 279648 416898
rect 310048 417454 310368 417486
rect 310048 417218 310090 417454
rect 310326 417218 310368 417454
rect 310048 417134 310368 417218
rect 310048 416898 310090 417134
rect 310326 416898 310368 417134
rect 310048 416866 310368 416898
rect 340768 417454 341088 417486
rect 340768 417218 340810 417454
rect 341046 417218 341088 417454
rect 340768 417134 341088 417218
rect 340768 416898 340810 417134
rect 341046 416898 341088 417134
rect 340768 416866 341088 416898
rect 371488 417454 371808 417486
rect 371488 417218 371530 417454
rect 371766 417218 371808 417454
rect 371488 417134 371808 417218
rect 371488 416898 371530 417134
rect 371766 416898 371808 417134
rect 371488 416866 371808 416898
rect 402208 417454 402528 417486
rect 402208 417218 402250 417454
rect 402486 417218 402528 417454
rect 402208 417134 402528 417218
rect 402208 416898 402250 417134
rect 402486 416898 402528 417134
rect 402208 416866 402528 416898
rect 432928 417454 433248 417486
rect 432928 417218 432970 417454
rect 433206 417218 433248 417454
rect 432928 417134 433248 417218
rect 432928 416898 432970 417134
rect 433206 416898 433248 417134
rect 432928 416866 433248 416898
rect 463648 417454 463968 417486
rect 463648 417218 463690 417454
rect 463926 417218 463968 417454
rect 463648 417134 463968 417218
rect 463648 416898 463690 417134
rect 463926 416898 463968 417134
rect 463648 416866 463968 416898
rect 494368 417454 494688 417486
rect 494368 417218 494410 417454
rect 494646 417218 494688 417454
rect 494368 417134 494688 417218
rect 494368 416898 494410 417134
rect 494646 416898 494688 417134
rect 494368 416866 494688 416898
rect 525088 417454 525408 417486
rect 525088 417218 525130 417454
rect 525366 417218 525408 417454
rect 525088 417134 525408 417218
rect 525088 416898 525130 417134
rect 525366 416898 525408 417134
rect 525088 416866 525408 416898
rect 48928 399454 49248 399486
rect 48928 399218 48970 399454
rect 49206 399218 49248 399454
rect 48928 399134 49248 399218
rect 48928 398898 48970 399134
rect 49206 398898 49248 399134
rect 48928 398866 49248 398898
rect 79648 399454 79968 399486
rect 79648 399218 79690 399454
rect 79926 399218 79968 399454
rect 79648 399134 79968 399218
rect 79648 398898 79690 399134
rect 79926 398898 79968 399134
rect 79648 398866 79968 398898
rect 110368 399454 110688 399486
rect 110368 399218 110410 399454
rect 110646 399218 110688 399454
rect 110368 399134 110688 399218
rect 110368 398898 110410 399134
rect 110646 398898 110688 399134
rect 110368 398866 110688 398898
rect 141088 399454 141408 399486
rect 141088 399218 141130 399454
rect 141366 399218 141408 399454
rect 141088 399134 141408 399218
rect 141088 398898 141130 399134
rect 141366 398898 141408 399134
rect 141088 398866 141408 398898
rect 171808 399454 172128 399486
rect 171808 399218 171850 399454
rect 172086 399218 172128 399454
rect 171808 399134 172128 399218
rect 171808 398898 171850 399134
rect 172086 398898 172128 399134
rect 171808 398866 172128 398898
rect 202528 399454 202848 399486
rect 202528 399218 202570 399454
rect 202806 399218 202848 399454
rect 202528 399134 202848 399218
rect 202528 398898 202570 399134
rect 202806 398898 202848 399134
rect 202528 398866 202848 398898
rect 233248 399454 233568 399486
rect 233248 399218 233290 399454
rect 233526 399218 233568 399454
rect 233248 399134 233568 399218
rect 233248 398898 233290 399134
rect 233526 398898 233568 399134
rect 233248 398866 233568 398898
rect 263968 399454 264288 399486
rect 263968 399218 264010 399454
rect 264246 399218 264288 399454
rect 263968 399134 264288 399218
rect 263968 398898 264010 399134
rect 264246 398898 264288 399134
rect 263968 398866 264288 398898
rect 294688 399454 295008 399486
rect 294688 399218 294730 399454
rect 294966 399218 295008 399454
rect 294688 399134 295008 399218
rect 294688 398898 294730 399134
rect 294966 398898 295008 399134
rect 294688 398866 295008 398898
rect 325408 399454 325728 399486
rect 325408 399218 325450 399454
rect 325686 399218 325728 399454
rect 325408 399134 325728 399218
rect 325408 398898 325450 399134
rect 325686 398898 325728 399134
rect 325408 398866 325728 398898
rect 356128 399454 356448 399486
rect 356128 399218 356170 399454
rect 356406 399218 356448 399454
rect 356128 399134 356448 399218
rect 356128 398898 356170 399134
rect 356406 398898 356448 399134
rect 356128 398866 356448 398898
rect 386848 399454 387168 399486
rect 386848 399218 386890 399454
rect 387126 399218 387168 399454
rect 386848 399134 387168 399218
rect 386848 398898 386890 399134
rect 387126 398898 387168 399134
rect 386848 398866 387168 398898
rect 417568 399454 417888 399486
rect 417568 399218 417610 399454
rect 417846 399218 417888 399454
rect 417568 399134 417888 399218
rect 417568 398898 417610 399134
rect 417846 398898 417888 399134
rect 417568 398866 417888 398898
rect 448288 399454 448608 399486
rect 448288 399218 448330 399454
rect 448566 399218 448608 399454
rect 448288 399134 448608 399218
rect 448288 398898 448330 399134
rect 448566 398898 448608 399134
rect 448288 398866 448608 398898
rect 479008 399454 479328 399486
rect 479008 399218 479050 399454
rect 479286 399218 479328 399454
rect 479008 399134 479328 399218
rect 479008 398898 479050 399134
rect 479286 398898 479328 399134
rect 479008 398866 479328 398898
rect 509728 399454 510048 399486
rect 509728 399218 509770 399454
rect 510006 399218 510048 399454
rect 509728 399134 510048 399218
rect 509728 398898 509770 399134
rect 510006 398898 510048 399134
rect 509728 398866 510048 398898
rect 33568 381454 33888 381486
rect 33568 381218 33610 381454
rect 33846 381218 33888 381454
rect 33568 381134 33888 381218
rect 33568 380898 33610 381134
rect 33846 380898 33888 381134
rect 33568 380866 33888 380898
rect 64288 381454 64608 381486
rect 64288 381218 64330 381454
rect 64566 381218 64608 381454
rect 64288 381134 64608 381218
rect 64288 380898 64330 381134
rect 64566 380898 64608 381134
rect 64288 380866 64608 380898
rect 95008 381454 95328 381486
rect 95008 381218 95050 381454
rect 95286 381218 95328 381454
rect 95008 381134 95328 381218
rect 95008 380898 95050 381134
rect 95286 380898 95328 381134
rect 95008 380866 95328 380898
rect 125728 381454 126048 381486
rect 125728 381218 125770 381454
rect 126006 381218 126048 381454
rect 125728 381134 126048 381218
rect 125728 380898 125770 381134
rect 126006 380898 126048 381134
rect 125728 380866 126048 380898
rect 156448 381454 156768 381486
rect 156448 381218 156490 381454
rect 156726 381218 156768 381454
rect 156448 381134 156768 381218
rect 156448 380898 156490 381134
rect 156726 380898 156768 381134
rect 156448 380866 156768 380898
rect 187168 381454 187488 381486
rect 187168 381218 187210 381454
rect 187446 381218 187488 381454
rect 187168 381134 187488 381218
rect 187168 380898 187210 381134
rect 187446 380898 187488 381134
rect 187168 380866 187488 380898
rect 217888 381454 218208 381486
rect 217888 381218 217930 381454
rect 218166 381218 218208 381454
rect 217888 381134 218208 381218
rect 217888 380898 217930 381134
rect 218166 380898 218208 381134
rect 217888 380866 218208 380898
rect 248608 381454 248928 381486
rect 248608 381218 248650 381454
rect 248886 381218 248928 381454
rect 248608 381134 248928 381218
rect 248608 380898 248650 381134
rect 248886 380898 248928 381134
rect 248608 380866 248928 380898
rect 279328 381454 279648 381486
rect 279328 381218 279370 381454
rect 279606 381218 279648 381454
rect 279328 381134 279648 381218
rect 279328 380898 279370 381134
rect 279606 380898 279648 381134
rect 279328 380866 279648 380898
rect 310048 381454 310368 381486
rect 310048 381218 310090 381454
rect 310326 381218 310368 381454
rect 310048 381134 310368 381218
rect 310048 380898 310090 381134
rect 310326 380898 310368 381134
rect 310048 380866 310368 380898
rect 340768 381454 341088 381486
rect 340768 381218 340810 381454
rect 341046 381218 341088 381454
rect 340768 381134 341088 381218
rect 340768 380898 340810 381134
rect 341046 380898 341088 381134
rect 340768 380866 341088 380898
rect 371488 381454 371808 381486
rect 371488 381218 371530 381454
rect 371766 381218 371808 381454
rect 371488 381134 371808 381218
rect 371488 380898 371530 381134
rect 371766 380898 371808 381134
rect 371488 380866 371808 380898
rect 402208 381454 402528 381486
rect 402208 381218 402250 381454
rect 402486 381218 402528 381454
rect 402208 381134 402528 381218
rect 402208 380898 402250 381134
rect 402486 380898 402528 381134
rect 402208 380866 402528 380898
rect 432928 381454 433248 381486
rect 432928 381218 432970 381454
rect 433206 381218 433248 381454
rect 432928 381134 433248 381218
rect 432928 380898 432970 381134
rect 433206 380898 433248 381134
rect 432928 380866 433248 380898
rect 463648 381454 463968 381486
rect 463648 381218 463690 381454
rect 463926 381218 463968 381454
rect 463648 381134 463968 381218
rect 463648 380898 463690 381134
rect 463926 380898 463968 381134
rect 463648 380866 463968 380898
rect 494368 381454 494688 381486
rect 494368 381218 494410 381454
rect 494646 381218 494688 381454
rect 494368 381134 494688 381218
rect 494368 380898 494410 381134
rect 494646 380898 494688 381134
rect 494368 380866 494688 380898
rect 525088 381454 525408 381486
rect 525088 381218 525130 381454
rect 525366 381218 525408 381454
rect 525088 381134 525408 381218
rect 525088 380898 525130 381134
rect 525366 380898 525408 381134
rect 525088 380866 525408 380898
rect 48928 363454 49248 363486
rect 48928 363218 48970 363454
rect 49206 363218 49248 363454
rect 48928 363134 49248 363218
rect 48928 362898 48970 363134
rect 49206 362898 49248 363134
rect 48928 362866 49248 362898
rect 79648 363454 79968 363486
rect 79648 363218 79690 363454
rect 79926 363218 79968 363454
rect 79648 363134 79968 363218
rect 79648 362898 79690 363134
rect 79926 362898 79968 363134
rect 79648 362866 79968 362898
rect 110368 363454 110688 363486
rect 110368 363218 110410 363454
rect 110646 363218 110688 363454
rect 110368 363134 110688 363218
rect 110368 362898 110410 363134
rect 110646 362898 110688 363134
rect 110368 362866 110688 362898
rect 141088 363454 141408 363486
rect 141088 363218 141130 363454
rect 141366 363218 141408 363454
rect 141088 363134 141408 363218
rect 141088 362898 141130 363134
rect 141366 362898 141408 363134
rect 141088 362866 141408 362898
rect 171808 363454 172128 363486
rect 171808 363218 171850 363454
rect 172086 363218 172128 363454
rect 171808 363134 172128 363218
rect 171808 362898 171850 363134
rect 172086 362898 172128 363134
rect 171808 362866 172128 362898
rect 202528 363454 202848 363486
rect 202528 363218 202570 363454
rect 202806 363218 202848 363454
rect 202528 363134 202848 363218
rect 202528 362898 202570 363134
rect 202806 362898 202848 363134
rect 202528 362866 202848 362898
rect 233248 363454 233568 363486
rect 233248 363218 233290 363454
rect 233526 363218 233568 363454
rect 233248 363134 233568 363218
rect 233248 362898 233290 363134
rect 233526 362898 233568 363134
rect 233248 362866 233568 362898
rect 263968 363454 264288 363486
rect 263968 363218 264010 363454
rect 264246 363218 264288 363454
rect 263968 363134 264288 363218
rect 263968 362898 264010 363134
rect 264246 362898 264288 363134
rect 263968 362866 264288 362898
rect 294688 363454 295008 363486
rect 294688 363218 294730 363454
rect 294966 363218 295008 363454
rect 294688 363134 295008 363218
rect 294688 362898 294730 363134
rect 294966 362898 295008 363134
rect 294688 362866 295008 362898
rect 325408 363454 325728 363486
rect 325408 363218 325450 363454
rect 325686 363218 325728 363454
rect 325408 363134 325728 363218
rect 325408 362898 325450 363134
rect 325686 362898 325728 363134
rect 325408 362866 325728 362898
rect 356128 363454 356448 363486
rect 356128 363218 356170 363454
rect 356406 363218 356448 363454
rect 356128 363134 356448 363218
rect 356128 362898 356170 363134
rect 356406 362898 356448 363134
rect 356128 362866 356448 362898
rect 386848 363454 387168 363486
rect 386848 363218 386890 363454
rect 387126 363218 387168 363454
rect 386848 363134 387168 363218
rect 386848 362898 386890 363134
rect 387126 362898 387168 363134
rect 386848 362866 387168 362898
rect 417568 363454 417888 363486
rect 417568 363218 417610 363454
rect 417846 363218 417888 363454
rect 417568 363134 417888 363218
rect 417568 362898 417610 363134
rect 417846 362898 417888 363134
rect 417568 362866 417888 362898
rect 448288 363454 448608 363486
rect 448288 363218 448330 363454
rect 448566 363218 448608 363454
rect 448288 363134 448608 363218
rect 448288 362898 448330 363134
rect 448566 362898 448608 363134
rect 448288 362866 448608 362898
rect 479008 363454 479328 363486
rect 479008 363218 479050 363454
rect 479286 363218 479328 363454
rect 479008 363134 479328 363218
rect 479008 362898 479050 363134
rect 479286 362898 479328 363134
rect 479008 362866 479328 362898
rect 509728 363454 510048 363486
rect 509728 363218 509770 363454
rect 510006 363218 510048 363454
rect 509728 363134 510048 363218
rect 509728 362898 509770 363134
rect 510006 362898 510048 363134
rect 509728 362866 510048 362898
rect 33568 345454 33888 345486
rect 33568 345218 33610 345454
rect 33846 345218 33888 345454
rect 33568 345134 33888 345218
rect 33568 344898 33610 345134
rect 33846 344898 33888 345134
rect 33568 344866 33888 344898
rect 64288 345454 64608 345486
rect 64288 345218 64330 345454
rect 64566 345218 64608 345454
rect 64288 345134 64608 345218
rect 64288 344898 64330 345134
rect 64566 344898 64608 345134
rect 64288 344866 64608 344898
rect 95008 345454 95328 345486
rect 95008 345218 95050 345454
rect 95286 345218 95328 345454
rect 95008 345134 95328 345218
rect 95008 344898 95050 345134
rect 95286 344898 95328 345134
rect 95008 344866 95328 344898
rect 125728 345454 126048 345486
rect 125728 345218 125770 345454
rect 126006 345218 126048 345454
rect 125728 345134 126048 345218
rect 125728 344898 125770 345134
rect 126006 344898 126048 345134
rect 125728 344866 126048 344898
rect 156448 345454 156768 345486
rect 156448 345218 156490 345454
rect 156726 345218 156768 345454
rect 156448 345134 156768 345218
rect 156448 344898 156490 345134
rect 156726 344898 156768 345134
rect 156448 344866 156768 344898
rect 187168 345454 187488 345486
rect 187168 345218 187210 345454
rect 187446 345218 187488 345454
rect 187168 345134 187488 345218
rect 187168 344898 187210 345134
rect 187446 344898 187488 345134
rect 187168 344866 187488 344898
rect 217888 345454 218208 345486
rect 217888 345218 217930 345454
rect 218166 345218 218208 345454
rect 217888 345134 218208 345218
rect 217888 344898 217930 345134
rect 218166 344898 218208 345134
rect 217888 344866 218208 344898
rect 248608 345454 248928 345486
rect 248608 345218 248650 345454
rect 248886 345218 248928 345454
rect 248608 345134 248928 345218
rect 248608 344898 248650 345134
rect 248886 344898 248928 345134
rect 248608 344866 248928 344898
rect 279328 345454 279648 345486
rect 279328 345218 279370 345454
rect 279606 345218 279648 345454
rect 279328 345134 279648 345218
rect 279328 344898 279370 345134
rect 279606 344898 279648 345134
rect 279328 344866 279648 344898
rect 310048 345454 310368 345486
rect 310048 345218 310090 345454
rect 310326 345218 310368 345454
rect 310048 345134 310368 345218
rect 310048 344898 310090 345134
rect 310326 344898 310368 345134
rect 310048 344866 310368 344898
rect 340768 345454 341088 345486
rect 340768 345218 340810 345454
rect 341046 345218 341088 345454
rect 340768 345134 341088 345218
rect 340768 344898 340810 345134
rect 341046 344898 341088 345134
rect 340768 344866 341088 344898
rect 371488 345454 371808 345486
rect 371488 345218 371530 345454
rect 371766 345218 371808 345454
rect 371488 345134 371808 345218
rect 371488 344898 371530 345134
rect 371766 344898 371808 345134
rect 371488 344866 371808 344898
rect 402208 345454 402528 345486
rect 402208 345218 402250 345454
rect 402486 345218 402528 345454
rect 402208 345134 402528 345218
rect 402208 344898 402250 345134
rect 402486 344898 402528 345134
rect 402208 344866 402528 344898
rect 432928 345454 433248 345486
rect 432928 345218 432970 345454
rect 433206 345218 433248 345454
rect 432928 345134 433248 345218
rect 432928 344898 432970 345134
rect 433206 344898 433248 345134
rect 432928 344866 433248 344898
rect 463648 345454 463968 345486
rect 463648 345218 463690 345454
rect 463926 345218 463968 345454
rect 463648 345134 463968 345218
rect 463648 344898 463690 345134
rect 463926 344898 463968 345134
rect 463648 344866 463968 344898
rect 494368 345454 494688 345486
rect 494368 345218 494410 345454
rect 494646 345218 494688 345454
rect 494368 345134 494688 345218
rect 494368 344898 494410 345134
rect 494646 344898 494688 345134
rect 494368 344866 494688 344898
rect 525088 345454 525408 345486
rect 525088 345218 525130 345454
rect 525366 345218 525408 345454
rect 525088 345134 525408 345218
rect 525088 344898 525130 345134
rect 525366 344898 525408 345134
rect 525088 344866 525408 344898
rect 48928 327454 49248 327486
rect 48928 327218 48970 327454
rect 49206 327218 49248 327454
rect 48928 327134 49248 327218
rect 48928 326898 48970 327134
rect 49206 326898 49248 327134
rect 48928 326866 49248 326898
rect 79648 327454 79968 327486
rect 79648 327218 79690 327454
rect 79926 327218 79968 327454
rect 79648 327134 79968 327218
rect 79648 326898 79690 327134
rect 79926 326898 79968 327134
rect 79648 326866 79968 326898
rect 110368 327454 110688 327486
rect 110368 327218 110410 327454
rect 110646 327218 110688 327454
rect 110368 327134 110688 327218
rect 110368 326898 110410 327134
rect 110646 326898 110688 327134
rect 110368 326866 110688 326898
rect 141088 327454 141408 327486
rect 141088 327218 141130 327454
rect 141366 327218 141408 327454
rect 141088 327134 141408 327218
rect 141088 326898 141130 327134
rect 141366 326898 141408 327134
rect 141088 326866 141408 326898
rect 171808 327454 172128 327486
rect 171808 327218 171850 327454
rect 172086 327218 172128 327454
rect 171808 327134 172128 327218
rect 171808 326898 171850 327134
rect 172086 326898 172128 327134
rect 171808 326866 172128 326898
rect 202528 327454 202848 327486
rect 202528 327218 202570 327454
rect 202806 327218 202848 327454
rect 202528 327134 202848 327218
rect 202528 326898 202570 327134
rect 202806 326898 202848 327134
rect 202528 326866 202848 326898
rect 233248 327454 233568 327486
rect 233248 327218 233290 327454
rect 233526 327218 233568 327454
rect 233248 327134 233568 327218
rect 233248 326898 233290 327134
rect 233526 326898 233568 327134
rect 233248 326866 233568 326898
rect 263968 327454 264288 327486
rect 263968 327218 264010 327454
rect 264246 327218 264288 327454
rect 263968 327134 264288 327218
rect 263968 326898 264010 327134
rect 264246 326898 264288 327134
rect 263968 326866 264288 326898
rect 294688 327454 295008 327486
rect 294688 327218 294730 327454
rect 294966 327218 295008 327454
rect 294688 327134 295008 327218
rect 294688 326898 294730 327134
rect 294966 326898 295008 327134
rect 294688 326866 295008 326898
rect 325408 327454 325728 327486
rect 325408 327218 325450 327454
rect 325686 327218 325728 327454
rect 325408 327134 325728 327218
rect 325408 326898 325450 327134
rect 325686 326898 325728 327134
rect 325408 326866 325728 326898
rect 356128 327454 356448 327486
rect 356128 327218 356170 327454
rect 356406 327218 356448 327454
rect 356128 327134 356448 327218
rect 356128 326898 356170 327134
rect 356406 326898 356448 327134
rect 356128 326866 356448 326898
rect 386848 327454 387168 327486
rect 386848 327218 386890 327454
rect 387126 327218 387168 327454
rect 386848 327134 387168 327218
rect 386848 326898 386890 327134
rect 387126 326898 387168 327134
rect 386848 326866 387168 326898
rect 417568 327454 417888 327486
rect 417568 327218 417610 327454
rect 417846 327218 417888 327454
rect 417568 327134 417888 327218
rect 417568 326898 417610 327134
rect 417846 326898 417888 327134
rect 417568 326866 417888 326898
rect 448288 327454 448608 327486
rect 448288 327218 448330 327454
rect 448566 327218 448608 327454
rect 448288 327134 448608 327218
rect 448288 326898 448330 327134
rect 448566 326898 448608 327134
rect 448288 326866 448608 326898
rect 479008 327454 479328 327486
rect 479008 327218 479050 327454
rect 479286 327218 479328 327454
rect 479008 327134 479328 327218
rect 479008 326898 479050 327134
rect 479286 326898 479328 327134
rect 479008 326866 479328 326898
rect 509728 327454 510048 327486
rect 509728 327218 509770 327454
rect 510006 327218 510048 327454
rect 509728 327134 510048 327218
rect 509728 326898 509770 327134
rect 510006 326898 510048 327134
rect 509728 326866 510048 326898
rect 33568 309454 33888 309486
rect 33568 309218 33610 309454
rect 33846 309218 33888 309454
rect 33568 309134 33888 309218
rect 33568 308898 33610 309134
rect 33846 308898 33888 309134
rect 33568 308866 33888 308898
rect 64288 309454 64608 309486
rect 64288 309218 64330 309454
rect 64566 309218 64608 309454
rect 64288 309134 64608 309218
rect 64288 308898 64330 309134
rect 64566 308898 64608 309134
rect 64288 308866 64608 308898
rect 95008 309454 95328 309486
rect 95008 309218 95050 309454
rect 95286 309218 95328 309454
rect 95008 309134 95328 309218
rect 95008 308898 95050 309134
rect 95286 308898 95328 309134
rect 95008 308866 95328 308898
rect 125728 309454 126048 309486
rect 125728 309218 125770 309454
rect 126006 309218 126048 309454
rect 125728 309134 126048 309218
rect 125728 308898 125770 309134
rect 126006 308898 126048 309134
rect 125728 308866 126048 308898
rect 156448 309454 156768 309486
rect 156448 309218 156490 309454
rect 156726 309218 156768 309454
rect 156448 309134 156768 309218
rect 156448 308898 156490 309134
rect 156726 308898 156768 309134
rect 156448 308866 156768 308898
rect 187168 309454 187488 309486
rect 187168 309218 187210 309454
rect 187446 309218 187488 309454
rect 187168 309134 187488 309218
rect 187168 308898 187210 309134
rect 187446 308898 187488 309134
rect 187168 308866 187488 308898
rect 217888 309454 218208 309486
rect 217888 309218 217930 309454
rect 218166 309218 218208 309454
rect 217888 309134 218208 309218
rect 217888 308898 217930 309134
rect 218166 308898 218208 309134
rect 217888 308866 218208 308898
rect 248608 309454 248928 309486
rect 248608 309218 248650 309454
rect 248886 309218 248928 309454
rect 248608 309134 248928 309218
rect 248608 308898 248650 309134
rect 248886 308898 248928 309134
rect 248608 308866 248928 308898
rect 279328 309454 279648 309486
rect 279328 309218 279370 309454
rect 279606 309218 279648 309454
rect 279328 309134 279648 309218
rect 279328 308898 279370 309134
rect 279606 308898 279648 309134
rect 279328 308866 279648 308898
rect 310048 309454 310368 309486
rect 310048 309218 310090 309454
rect 310326 309218 310368 309454
rect 310048 309134 310368 309218
rect 310048 308898 310090 309134
rect 310326 308898 310368 309134
rect 310048 308866 310368 308898
rect 340768 309454 341088 309486
rect 340768 309218 340810 309454
rect 341046 309218 341088 309454
rect 340768 309134 341088 309218
rect 340768 308898 340810 309134
rect 341046 308898 341088 309134
rect 340768 308866 341088 308898
rect 371488 309454 371808 309486
rect 371488 309218 371530 309454
rect 371766 309218 371808 309454
rect 371488 309134 371808 309218
rect 371488 308898 371530 309134
rect 371766 308898 371808 309134
rect 371488 308866 371808 308898
rect 402208 309454 402528 309486
rect 402208 309218 402250 309454
rect 402486 309218 402528 309454
rect 402208 309134 402528 309218
rect 402208 308898 402250 309134
rect 402486 308898 402528 309134
rect 402208 308866 402528 308898
rect 432928 309454 433248 309486
rect 432928 309218 432970 309454
rect 433206 309218 433248 309454
rect 432928 309134 433248 309218
rect 432928 308898 432970 309134
rect 433206 308898 433248 309134
rect 432928 308866 433248 308898
rect 463648 309454 463968 309486
rect 463648 309218 463690 309454
rect 463926 309218 463968 309454
rect 463648 309134 463968 309218
rect 463648 308898 463690 309134
rect 463926 308898 463968 309134
rect 463648 308866 463968 308898
rect 494368 309454 494688 309486
rect 494368 309218 494410 309454
rect 494646 309218 494688 309454
rect 494368 309134 494688 309218
rect 494368 308898 494410 309134
rect 494646 308898 494688 309134
rect 494368 308866 494688 308898
rect 525088 309454 525408 309486
rect 525088 309218 525130 309454
rect 525366 309218 525408 309454
rect 525088 309134 525408 309218
rect 525088 308898 525130 309134
rect 525366 308898 525408 309134
rect 525088 308866 525408 308898
rect 48928 291454 49248 291486
rect 48928 291218 48970 291454
rect 49206 291218 49248 291454
rect 48928 291134 49248 291218
rect 48928 290898 48970 291134
rect 49206 290898 49248 291134
rect 48928 290866 49248 290898
rect 79648 291454 79968 291486
rect 79648 291218 79690 291454
rect 79926 291218 79968 291454
rect 79648 291134 79968 291218
rect 79648 290898 79690 291134
rect 79926 290898 79968 291134
rect 79648 290866 79968 290898
rect 110368 291454 110688 291486
rect 110368 291218 110410 291454
rect 110646 291218 110688 291454
rect 110368 291134 110688 291218
rect 110368 290898 110410 291134
rect 110646 290898 110688 291134
rect 110368 290866 110688 290898
rect 141088 291454 141408 291486
rect 141088 291218 141130 291454
rect 141366 291218 141408 291454
rect 141088 291134 141408 291218
rect 141088 290898 141130 291134
rect 141366 290898 141408 291134
rect 141088 290866 141408 290898
rect 171808 291454 172128 291486
rect 171808 291218 171850 291454
rect 172086 291218 172128 291454
rect 171808 291134 172128 291218
rect 171808 290898 171850 291134
rect 172086 290898 172128 291134
rect 171808 290866 172128 290898
rect 202528 291454 202848 291486
rect 202528 291218 202570 291454
rect 202806 291218 202848 291454
rect 202528 291134 202848 291218
rect 202528 290898 202570 291134
rect 202806 290898 202848 291134
rect 202528 290866 202848 290898
rect 233248 291454 233568 291486
rect 233248 291218 233290 291454
rect 233526 291218 233568 291454
rect 233248 291134 233568 291218
rect 233248 290898 233290 291134
rect 233526 290898 233568 291134
rect 233248 290866 233568 290898
rect 263968 291454 264288 291486
rect 263968 291218 264010 291454
rect 264246 291218 264288 291454
rect 263968 291134 264288 291218
rect 263968 290898 264010 291134
rect 264246 290898 264288 291134
rect 263968 290866 264288 290898
rect 294688 291454 295008 291486
rect 294688 291218 294730 291454
rect 294966 291218 295008 291454
rect 294688 291134 295008 291218
rect 294688 290898 294730 291134
rect 294966 290898 295008 291134
rect 294688 290866 295008 290898
rect 325408 291454 325728 291486
rect 325408 291218 325450 291454
rect 325686 291218 325728 291454
rect 325408 291134 325728 291218
rect 325408 290898 325450 291134
rect 325686 290898 325728 291134
rect 325408 290866 325728 290898
rect 356128 291454 356448 291486
rect 356128 291218 356170 291454
rect 356406 291218 356448 291454
rect 356128 291134 356448 291218
rect 356128 290898 356170 291134
rect 356406 290898 356448 291134
rect 356128 290866 356448 290898
rect 386848 291454 387168 291486
rect 386848 291218 386890 291454
rect 387126 291218 387168 291454
rect 386848 291134 387168 291218
rect 386848 290898 386890 291134
rect 387126 290898 387168 291134
rect 386848 290866 387168 290898
rect 417568 291454 417888 291486
rect 417568 291218 417610 291454
rect 417846 291218 417888 291454
rect 417568 291134 417888 291218
rect 417568 290898 417610 291134
rect 417846 290898 417888 291134
rect 417568 290866 417888 290898
rect 448288 291454 448608 291486
rect 448288 291218 448330 291454
rect 448566 291218 448608 291454
rect 448288 291134 448608 291218
rect 448288 290898 448330 291134
rect 448566 290898 448608 291134
rect 448288 290866 448608 290898
rect 479008 291454 479328 291486
rect 479008 291218 479050 291454
rect 479286 291218 479328 291454
rect 479008 291134 479328 291218
rect 479008 290898 479050 291134
rect 479286 290898 479328 291134
rect 479008 290866 479328 290898
rect 509728 291454 510048 291486
rect 509728 291218 509770 291454
rect 510006 291218 510048 291454
rect 509728 291134 510048 291218
rect 509728 290898 509770 291134
rect 510006 290898 510048 291134
rect 509728 290866 510048 290898
rect 33568 273454 33888 273486
rect 33568 273218 33610 273454
rect 33846 273218 33888 273454
rect 33568 273134 33888 273218
rect 33568 272898 33610 273134
rect 33846 272898 33888 273134
rect 33568 272866 33888 272898
rect 64288 273454 64608 273486
rect 64288 273218 64330 273454
rect 64566 273218 64608 273454
rect 64288 273134 64608 273218
rect 64288 272898 64330 273134
rect 64566 272898 64608 273134
rect 64288 272866 64608 272898
rect 95008 273454 95328 273486
rect 95008 273218 95050 273454
rect 95286 273218 95328 273454
rect 95008 273134 95328 273218
rect 95008 272898 95050 273134
rect 95286 272898 95328 273134
rect 95008 272866 95328 272898
rect 125728 273454 126048 273486
rect 125728 273218 125770 273454
rect 126006 273218 126048 273454
rect 125728 273134 126048 273218
rect 125728 272898 125770 273134
rect 126006 272898 126048 273134
rect 125728 272866 126048 272898
rect 156448 273454 156768 273486
rect 156448 273218 156490 273454
rect 156726 273218 156768 273454
rect 156448 273134 156768 273218
rect 156448 272898 156490 273134
rect 156726 272898 156768 273134
rect 156448 272866 156768 272898
rect 187168 273454 187488 273486
rect 187168 273218 187210 273454
rect 187446 273218 187488 273454
rect 187168 273134 187488 273218
rect 187168 272898 187210 273134
rect 187446 272898 187488 273134
rect 187168 272866 187488 272898
rect 217888 273454 218208 273486
rect 217888 273218 217930 273454
rect 218166 273218 218208 273454
rect 217888 273134 218208 273218
rect 217888 272898 217930 273134
rect 218166 272898 218208 273134
rect 217888 272866 218208 272898
rect 248608 273454 248928 273486
rect 248608 273218 248650 273454
rect 248886 273218 248928 273454
rect 248608 273134 248928 273218
rect 248608 272898 248650 273134
rect 248886 272898 248928 273134
rect 248608 272866 248928 272898
rect 279328 273454 279648 273486
rect 279328 273218 279370 273454
rect 279606 273218 279648 273454
rect 279328 273134 279648 273218
rect 279328 272898 279370 273134
rect 279606 272898 279648 273134
rect 279328 272866 279648 272898
rect 310048 273454 310368 273486
rect 310048 273218 310090 273454
rect 310326 273218 310368 273454
rect 310048 273134 310368 273218
rect 310048 272898 310090 273134
rect 310326 272898 310368 273134
rect 310048 272866 310368 272898
rect 340768 273454 341088 273486
rect 340768 273218 340810 273454
rect 341046 273218 341088 273454
rect 340768 273134 341088 273218
rect 340768 272898 340810 273134
rect 341046 272898 341088 273134
rect 340768 272866 341088 272898
rect 371488 273454 371808 273486
rect 371488 273218 371530 273454
rect 371766 273218 371808 273454
rect 371488 273134 371808 273218
rect 371488 272898 371530 273134
rect 371766 272898 371808 273134
rect 371488 272866 371808 272898
rect 402208 273454 402528 273486
rect 402208 273218 402250 273454
rect 402486 273218 402528 273454
rect 402208 273134 402528 273218
rect 402208 272898 402250 273134
rect 402486 272898 402528 273134
rect 402208 272866 402528 272898
rect 432928 273454 433248 273486
rect 432928 273218 432970 273454
rect 433206 273218 433248 273454
rect 432928 273134 433248 273218
rect 432928 272898 432970 273134
rect 433206 272898 433248 273134
rect 432928 272866 433248 272898
rect 463648 273454 463968 273486
rect 463648 273218 463690 273454
rect 463926 273218 463968 273454
rect 463648 273134 463968 273218
rect 463648 272898 463690 273134
rect 463926 272898 463968 273134
rect 463648 272866 463968 272898
rect 494368 273454 494688 273486
rect 494368 273218 494410 273454
rect 494646 273218 494688 273454
rect 494368 273134 494688 273218
rect 494368 272898 494410 273134
rect 494646 272898 494688 273134
rect 494368 272866 494688 272898
rect 525088 273454 525408 273486
rect 525088 273218 525130 273454
rect 525366 273218 525408 273454
rect 525088 273134 525408 273218
rect 525088 272898 525130 273134
rect 525366 272898 525408 273134
rect 525088 272866 525408 272898
rect 48928 255454 49248 255486
rect 48928 255218 48970 255454
rect 49206 255218 49248 255454
rect 48928 255134 49248 255218
rect 48928 254898 48970 255134
rect 49206 254898 49248 255134
rect 48928 254866 49248 254898
rect 79648 255454 79968 255486
rect 79648 255218 79690 255454
rect 79926 255218 79968 255454
rect 79648 255134 79968 255218
rect 79648 254898 79690 255134
rect 79926 254898 79968 255134
rect 79648 254866 79968 254898
rect 110368 255454 110688 255486
rect 110368 255218 110410 255454
rect 110646 255218 110688 255454
rect 110368 255134 110688 255218
rect 110368 254898 110410 255134
rect 110646 254898 110688 255134
rect 110368 254866 110688 254898
rect 141088 255454 141408 255486
rect 141088 255218 141130 255454
rect 141366 255218 141408 255454
rect 141088 255134 141408 255218
rect 141088 254898 141130 255134
rect 141366 254898 141408 255134
rect 141088 254866 141408 254898
rect 171808 255454 172128 255486
rect 171808 255218 171850 255454
rect 172086 255218 172128 255454
rect 171808 255134 172128 255218
rect 171808 254898 171850 255134
rect 172086 254898 172128 255134
rect 171808 254866 172128 254898
rect 202528 255454 202848 255486
rect 202528 255218 202570 255454
rect 202806 255218 202848 255454
rect 202528 255134 202848 255218
rect 202528 254898 202570 255134
rect 202806 254898 202848 255134
rect 202528 254866 202848 254898
rect 233248 255454 233568 255486
rect 233248 255218 233290 255454
rect 233526 255218 233568 255454
rect 233248 255134 233568 255218
rect 233248 254898 233290 255134
rect 233526 254898 233568 255134
rect 233248 254866 233568 254898
rect 263968 255454 264288 255486
rect 263968 255218 264010 255454
rect 264246 255218 264288 255454
rect 263968 255134 264288 255218
rect 263968 254898 264010 255134
rect 264246 254898 264288 255134
rect 263968 254866 264288 254898
rect 294688 255454 295008 255486
rect 294688 255218 294730 255454
rect 294966 255218 295008 255454
rect 294688 255134 295008 255218
rect 294688 254898 294730 255134
rect 294966 254898 295008 255134
rect 294688 254866 295008 254898
rect 325408 255454 325728 255486
rect 325408 255218 325450 255454
rect 325686 255218 325728 255454
rect 325408 255134 325728 255218
rect 325408 254898 325450 255134
rect 325686 254898 325728 255134
rect 325408 254866 325728 254898
rect 356128 255454 356448 255486
rect 356128 255218 356170 255454
rect 356406 255218 356448 255454
rect 356128 255134 356448 255218
rect 356128 254898 356170 255134
rect 356406 254898 356448 255134
rect 356128 254866 356448 254898
rect 386848 255454 387168 255486
rect 386848 255218 386890 255454
rect 387126 255218 387168 255454
rect 386848 255134 387168 255218
rect 386848 254898 386890 255134
rect 387126 254898 387168 255134
rect 386848 254866 387168 254898
rect 417568 255454 417888 255486
rect 417568 255218 417610 255454
rect 417846 255218 417888 255454
rect 417568 255134 417888 255218
rect 417568 254898 417610 255134
rect 417846 254898 417888 255134
rect 417568 254866 417888 254898
rect 448288 255454 448608 255486
rect 448288 255218 448330 255454
rect 448566 255218 448608 255454
rect 448288 255134 448608 255218
rect 448288 254898 448330 255134
rect 448566 254898 448608 255134
rect 448288 254866 448608 254898
rect 479008 255454 479328 255486
rect 479008 255218 479050 255454
rect 479286 255218 479328 255454
rect 479008 255134 479328 255218
rect 479008 254898 479050 255134
rect 479286 254898 479328 255134
rect 479008 254866 479328 254898
rect 509728 255454 510048 255486
rect 509728 255218 509770 255454
rect 510006 255218 510048 255454
rect 509728 255134 510048 255218
rect 509728 254898 509770 255134
rect 510006 254898 510048 255134
rect 509728 254866 510048 254898
rect 33568 237454 33888 237486
rect 33568 237218 33610 237454
rect 33846 237218 33888 237454
rect 33568 237134 33888 237218
rect 33568 236898 33610 237134
rect 33846 236898 33888 237134
rect 33568 236866 33888 236898
rect 64288 237454 64608 237486
rect 64288 237218 64330 237454
rect 64566 237218 64608 237454
rect 64288 237134 64608 237218
rect 64288 236898 64330 237134
rect 64566 236898 64608 237134
rect 64288 236866 64608 236898
rect 95008 237454 95328 237486
rect 95008 237218 95050 237454
rect 95286 237218 95328 237454
rect 95008 237134 95328 237218
rect 95008 236898 95050 237134
rect 95286 236898 95328 237134
rect 95008 236866 95328 236898
rect 125728 237454 126048 237486
rect 125728 237218 125770 237454
rect 126006 237218 126048 237454
rect 125728 237134 126048 237218
rect 125728 236898 125770 237134
rect 126006 236898 126048 237134
rect 125728 236866 126048 236898
rect 156448 237454 156768 237486
rect 156448 237218 156490 237454
rect 156726 237218 156768 237454
rect 156448 237134 156768 237218
rect 156448 236898 156490 237134
rect 156726 236898 156768 237134
rect 156448 236866 156768 236898
rect 187168 237454 187488 237486
rect 187168 237218 187210 237454
rect 187446 237218 187488 237454
rect 187168 237134 187488 237218
rect 187168 236898 187210 237134
rect 187446 236898 187488 237134
rect 187168 236866 187488 236898
rect 217888 237454 218208 237486
rect 217888 237218 217930 237454
rect 218166 237218 218208 237454
rect 217888 237134 218208 237218
rect 217888 236898 217930 237134
rect 218166 236898 218208 237134
rect 217888 236866 218208 236898
rect 248608 237454 248928 237486
rect 248608 237218 248650 237454
rect 248886 237218 248928 237454
rect 248608 237134 248928 237218
rect 248608 236898 248650 237134
rect 248886 236898 248928 237134
rect 248608 236866 248928 236898
rect 279328 237454 279648 237486
rect 279328 237218 279370 237454
rect 279606 237218 279648 237454
rect 279328 237134 279648 237218
rect 279328 236898 279370 237134
rect 279606 236898 279648 237134
rect 279328 236866 279648 236898
rect 310048 237454 310368 237486
rect 310048 237218 310090 237454
rect 310326 237218 310368 237454
rect 310048 237134 310368 237218
rect 310048 236898 310090 237134
rect 310326 236898 310368 237134
rect 310048 236866 310368 236898
rect 340768 237454 341088 237486
rect 340768 237218 340810 237454
rect 341046 237218 341088 237454
rect 340768 237134 341088 237218
rect 340768 236898 340810 237134
rect 341046 236898 341088 237134
rect 340768 236866 341088 236898
rect 371488 237454 371808 237486
rect 371488 237218 371530 237454
rect 371766 237218 371808 237454
rect 371488 237134 371808 237218
rect 371488 236898 371530 237134
rect 371766 236898 371808 237134
rect 371488 236866 371808 236898
rect 402208 237454 402528 237486
rect 402208 237218 402250 237454
rect 402486 237218 402528 237454
rect 402208 237134 402528 237218
rect 402208 236898 402250 237134
rect 402486 236898 402528 237134
rect 402208 236866 402528 236898
rect 432928 237454 433248 237486
rect 432928 237218 432970 237454
rect 433206 237218 433248 237454
rect 432928 237134 433248 237218
rect 432928 236898 432970 237134
rect 433206 236898 433248 237134
rect 432928 236866 433248 236898
rect 463648 237454 463968 237486
rect 463648 237218 463690 237454
rect 463926 237218 463968 237454
rect 463648 237134 463968 237218
rect 463648 236898 463690 237134
rect 463926 236898 463968 237134
rect 463648 236866 463968 236898
rect 494368 237454 494688 237486
rect 494368 237218 494410 237454
rect 494646 237218 494688 237454
rect 494368 237134 494688 237218
rect 494368 236898 494410 237134
rect 494646 236898 494688 237134
rect 494368 236866 494688 236898
rect 525088 237454 525408 237486
rect 525088 237218 525130 237454
rect 525366 237218 525408 237454
rect 525088 237134 525408 237218
rect 525088 236898 525130 237134
rect 525366 236898 525408 237134
rect 525088 236866 525408 236898
rect 48928 219454 49248 219486
rect 48928 219218 48970 219454
rect 49206 219218 49248 219454
rect 48928 219134 49248 219218
rect 48928 218898 48970 219134
rect 49206 218898 49248 219134
rect 48928 218866 49248 218898
rect 79648 219454 79968 219486
rect 79648 219218 79690 219454
rect 79926 219218 79968 219454
rect 79648 219134 79968 219218
rect 79648 218898 79690 219134
rect 79926 218898 79968 219134
rect 79648 218866 79968 218898
rect 110368 219454 110688 219486
rect 110368 219218 110410 219454
rect 110646 219218 110688 219454
rect 110368 219134 110688 219218
rect 110368 218898 110410 219134
rect 110646 218898 110688 219134
rect 110368 218866 110688 218898
rect 141088 219454 141408 219486
rect 141088 219218 141130 219454
rect 141366 219218 141408 219454
rect 141088 219134 141408 219218
rect 141088 218898 141130 219134
rect 141366 218898 141408 219134
rect 141088 218866 141408 218898
rect 171808 219454 172128 219486
rect 171808 219218 171850 219454
rect 172086 219218 172128 219454
rect 171808 219134 172128 219218
rect 171808 218898 171850 219134
rect 172086 218898 172128 219134
rect 171808 218866 172128 218898
rect 202528 219454 202848 219486
rect 202528 219218 202570 219454
rect 202806 219218 202848 219454
rect 202528 219134 202848 219218
rect 202528 218898 202570 219134
rect 202806 218898 202848 219134
rect 202528 218866 202848 218898
rect 233248 219454 233568 219486
rect 233248 219218 233290 219454
rect 233526 219218 233568 219454
rect 233248 219134 233568 219218
rect 233248 218898 233290 219134
rect 233526 218898 233568 219134
rect 233248 218866 233568 218898
rect 263968 219454 264288 219486
rect 263968 219218 264010 219454
rect 264246 219218 264288 219454
rect 263968 219134 264288 219218
rect 263968 218898 264010 219134
rect 264246 218898 264288 219134
rect 263968 218866 264288 218898
rect 294688 219454 295008 219486
rect 294688 219218 294730 219454
rect 294966 219218 295008 219454
rect 294688 219134 295008 219218
rect 294688 218898 294730 219134
rect 294966 218898 295008 219134
rect 294688 218866 295008 218898
rect 325408 219454 325728 219486
rect 325408 219218 325450 219454
rect 325686 219218 325728 219454
rect 325408 219134 325728 219218
rect 325408 218898 325450 219134
rect 325686 218898 325728 219134
rect 325408 218866 325728 218898
rect 356128 219454 356448 219486
rect 356128 219218 356170 219454
rect 356406 219218 356448 219454
rect 356128 219134 356448 219218
rect 356128 218898 356170 219134
rect 356406 218898 356448 219134
rect 356128 218866 356448 218898
rect 386848 219454 387168 219486
rect 386848 219218 386890 219454
rect 387126 219218 387168 219454
rect 386848 219134 387168 219218
rect 386848 218898 386890 219134
rect 387126 218898 387168 219134
rect 386848 218866 387168 218898
rect 417568 219454 417888 219486
rect 417568 219218 417610 219454
rect 417846 219218 417888 219454
rect 417568 219134 417888 219218
rect 417568 218898 417610 219134
rect 417846 218898 417888 219134
rect 417568 218866 417888 218898
rect 448288 219454 448608 219486
rect 448288 219218 448330 219454
rect 448566 219218 448608 219454
rect 448288 219134 448608 219218
rect 448288 218898 448330 219134
rect 448566 218898 448608 219134
rect 448288 218866 448608 218898
rect 479008 219454 479328 219486
rect 479008 219218 479050 219454
rect 479286 219218 479328 219454
rect 479008 219134 479328 219218
rect 479008 218898 479050 219134
rect 479286 218898 479328 219134
rect 479008 218866 479328 218898
rect 509728 219454 510048 219486
rect 509728 219218 509770 219454
rect 510006 219218 510048 219454
rect 509728 219134 510048 219218
rect 509728 218898 509770 219134
rect 510006 218898 510048 219134
rect 509728 218866 510048 218898
rect 33568 201454 33888 201486
rect 33568 201218 33610 201454
rect 33846 201218 33888 201454
rect 33568 201134 33888 201218
rect 33568 200898 33610 201134
rect 33846 200898 33888 201134
rect 33568 200866 33888 200898
rect 64288 201454 64608 201486
rect 64288 201218 64330 201454
rect 64566 201218 64608 201454
rect 64288 201134 64608 201218
rect 64288 200898 64330 201134
rect 64566 200898 64608 201134
rect 64288 200866 64608 200898
rect 95008 201454 95328 201486
rect 95008 201218 95050 201454
rect 95286 201218 95328 201454
rect 95008 201134 95328 201218
rect 95008 200898 95050 201134
rect 95286 200898 95328 201134
rect 95008 200866 95328 200898
rect 125728 201454 126048 201486
rect 125728 201218 125770 201454
rect 126006 201218 126048 201454
rect 125728 201134 126048 201218
rect 125728 200898 125770 201134
rect 126006 200898 126048 201134
rect 125728 200866 126048 200898
rect 156448 201454 156768 201486
rect 156448 201218 156490 201454
rect 156726 201218 156768 201454
rect 156448 201134 156768 201218
rect 156448 200898 156490 201134
rect 156726 200898 156768 201134
rect 156448 200866 156768 200898
rect 187168 201454 187488 201486
rect 187168 201218 187210 201454
rect 187446 201218 187488 201454
rect 187168 201134 187488 201218
rect 187168 200898 187210 201134
rect 187446 200898 187488 201134
rect 187168 200866 187488 200898
rect 217888 201454 218208 201486
rect 217888 201218 217930 201454
rect 218166 201218 218208 201454
rect 217888 201134 218208 201218
rect 217888 200898 217930 201134
rect 218166 200898 218208 201134
rect 217888 200866 218208 200898
rect 248608 201454 248928 201486
rect 248608 201218 248650 201454
rect 248886 201218 248928 201454
rect 248608 201134 248928 201218
rect 248608 200898 248650 201134
rect 248886 200898 248928 201134
rect 248608 200866 248928 200898
rect 279328 201454 279648 201486
rect 279328 201218 279370 201454
rect 279606 201218 279648 201454
rect 279328 201134 279648 201218
rect 279328 200898 279370 201134
rect 279606 200898 279648 201134
rect 279328 200866 279648 200898
rect 310048 201454 310368 201486
rect 310048 201218 310090 201454
rect 310326 201218 310368 201454
rect 310048 201134 310368 201218
rect 310048 200898 310090 201134
rect 310326 200898 310368 201134
rect 310048 200866 310368 200898
rect 340768 201454 341088 201486
rect 340768 201218 340810 201454
rect 341046 201218 341088 201454
rect 340768 201134 341088 201218
rect 340768 200898 340810 201134
rect 341046 200898 341088 201134
rect 340768 200866 341088 200898
rect 371488 201454 371808 201486
rect 371488 201218 371530 201454
rect 371766 201218 371808 201454
rect 371488 201134 371808 201218
rect 371488 200898 371530 201134
rect 371766 200898 371808 201134
rect 371488 200866 371808 200898
rect 402208 201454 402528 201486
rect 402208 201218 402250 201454
rect 402486 201218 402528 201454
rect 402208 201134 402528 201218
rect 402208 200898 402250 201134
rect 402486 200898 402528 201134
rect 402208 200866 402528 200898
rect 432928 201454 433248 201486
rect 432928 201218 432970 201454
rect 433206 201218 433248 201454
rect 432928 201134 433248 201218
rect 432928 200898 432970 201134
rect 433206 200898 433248 201134
rect 432928 200866 433248 200898
rect 463648 201454 463968 201486
rect 463648 201218 463690 201454
rect 463926 201218 463968 201454
rect 463648 201134 463968 201218
rect 463648 200898 463690 201134
rect 463926 200898 463968 201134
rect 463648 200866 463968 200898
rect 494368 201454 494688 201486
rect 494368 201218 494410 201454
rect 494646 201218 494688 201454
rect 494368 201134 494688 201218
rect 494368 200898 494410 201134
rect 494646 200898 494688 201134
rect 494368 200866 494688 200898
rect 525088 201454 525408 201486
rect 525088 201218 525130 201454
rect 525366 201218 525408 201454
rect 525088 201134 525408 201218
rect 525088 200898 525130 201134
rect 525366 200898 525408 201134
rect 525088 200866 525408 200898
rect 48928 183454 49248 183486
rect 48928 183218 48970 183454
rect 49206 183218 49248 183454
rect 48928 183134 49248 183218
rect 48928 182898 48970 183134
rect 49206 182898 49248 183134
rect 48928 182866 49248 182898
rect 79648 183454 79968 183486
rect 79648 183218 79690 183454
rect 79926 183218 79968 183454
rect 79648 183134 79968 183218
rect 79648 182898 79690 183134
rect 79926 182898 79968 183134
rect 79648 182866 79968 182898
rect 110368 183454 110688 183486
rect 110368 183218 110410 183454
rect 110646 183218 110688 183454
rect 110368 183134 110688 183218
rect 110368 182898 110410 183134
rect 110646 182898 110688 183134
rect 110368 182866 110688 182898
rect 141088 183454 141408 183486
rect 141088 183218 141130 183454
rect 141366 183218 141408 183454
rect 141088 183134 141408 183218
rect 141088 182898 141130 183134
rect 141366 182898 141408 183134
rect 141088 182866 141408 182898
rect 171808 183454 172128 183486
rect 171808 183218 171850 183454
rect 172086 183218 172128 183454
rect 171808 183134 172128 183218
rect 171808 182898 171850 183134
rect 172086 182898 172128 183134
rect 171808 182866 172128 182898
rect 202528 183454 202848 183486
rect 202528 183218 202570 183454
rect 202806 183218 202848 183454
rect 202528 183134 202848 183218
rect 202528 182898 202570 183134
rect 202806 182898 202848 183134
rect 202528 182866 202848 182898
rect 233248 183454 233568 183486
rect 233248 183218 233290 183454
rect 233526 183218 233568 183454
rect 233248 183134 233568 183218
rect 233248 182898 233290 183134
rect 233526 182898 233568 183134
rect 233248 182866 233568 182898
rect 263968 183454 264288 183486
rect 263968 183218 264010 183454
rect 264246 183218 264288 183454
rect 263968 183134 264288 183218
rect 263968 182898 264010 183134
rect 264246 182898 264288 183134
rect 263968 182866 264288 182898
rect 294688 183454 295008 183486
rect 294688 183218 294730 183454
rect 294966 183218 295008 183454
rect 294688 183134 295008 183218
rect 294688 182898 294730 183134
rect 294966 182898 295008 183134
rect 294688 182866 295008 182898
rect 325408 183454 325728 183486
rect 325408 183218 325450 183454
rect 325686 183218 325728 183454
rect 325408 183134 325728 183218
rect 325408 182898 325450 183134
rect 325686 182898 325728 183134
rect 325408 182866 325728 182898
rect 356128 183454 356448 183486
rect 356128 183218 356170 183454
rect 356406 183218 356448 183454
rect 356128 183134 356448 183218
rect 356128 182898 356170 183134
rect 356406 182898 356448 183134
rect 356128 182866 356448 182898
rect 386848 183454 387168 183486
rect 386848 183218 386890 183454
rect 387126 183218 387168 183454
rect 386848 183134 387168 183218
rect 386848 182898 386890 183134
rect 387126 182898 387168 183134
rect 386848 182866 387168 182898
rect 417568 183454 417888 183486
rect 417568 183218 417610 183454
rect 417846 183218 417888 183454
rect 417568 183134 417888 183218
rect 417568 182898 417610 183134
rect 417846 182898 417888 183134
rect 417568 182866 417888 182898
rect 448288 183454 448608 183486
rect 448288 183218 448330 183454
rect 448566 183218 448608 183454
rect 448288 183134 448608 183218
rect 448288 182898 448330 183134
rect 448566 182898 448608 183134
rect 448288 182866 448608 182898
rect 479008 183454 479328 183486
rect 479008 183218 479050 183454
rect 479286 183218 479328 183454
rect 479008 183134 479328 183218
rect 479008 182898 479050 183134
rect 479286 182898 479328 183134
rect 479008 182866 479328 182898
rect 509728 183454 510048 183486
rect 509728 183218 509770 183454
rect 510006 183218 510048 183454
rect 509728 183134 510048 183218
rect 509728 182898 509770 183134
rect 510006 182898 510048 183134
rect 509728 182866 510048 182898
rect 33568 165454 33888 165486
rect 33568 165218 33610 165454
rect 33846 165218 33888 165454
rect 33568 165134 33888 165218
rect 33568 164898 33610 165134
rect 33846 164898 33888 165134
rect 33568 164866 33888 164898
rect 64288 165454 64608 165486
rect 64288 165218 64330 165454
rect 64566 165218 64608 165454
rect 64288 165134 64608 165218
rect 64288 164898 64330 165134
rect 64566 164898 64608 165134
rect 64288 164866 64608 164898
rect 95008 165454 95328 165486
rect 95008 165218 95050 165454
rect 95286 165218 95328 165454
rect 95008 165134 95328 165218
rect 95008 164898 95050 165134
rect 95286 164898 95328 165134
rect 95008 164866 95328 164898
rect 125728 165454 126048 165486
rect 125728 165218 125770 165454
rect 126006 165218 126048 165454
rect 125728 165134 126048 165218
rect 125728 164898 125770 165134
rect 126006 164898 126048 165134
rect 125728 164866 126048 164898
rect 156448 165454 156768 165486
rect 156448 165218 156490 165454
rect 156726 165218 156768 165454
rect 156448 165134 156768 165218
rect 156448 164898 156490 165134
rect 156726 164898 156768 165134
rect 156448 164866 156768 164898
rect 187168 165454 187488 165486
rect 187168 165218 187210 165454
rect 187446 165218 187488 165454
rect 187168 165134 187488 165218
rect 187168 164898 187210 165134
rect 187446 164898 187488 165134
rect 187168 164866 187488 164898
rect 217888 165454 218208 165486
rect 217888 165218 217930 165454
rect 218166 165218 218208 165454
rect 217888 165134 218208 165218
rect 217888 164898 217930 165134
rect 218166 164898 218208 165134
rect 217888 164866 218208 164898
rect 248608 165454 248928 165486
rect 248608 165218 248650 165454
rect 248886 165218 248928 165454
rect 248608 165134 248928 165218
rect 248608 164898 248650 165134
rect 248886 164898 248928 165134
rect 248608 164866 248928 164898
rect 279328 165454 279648 165486
rect 279328 165218 279370 165454
rect 279606 165218 279648 165454
rect 279328 165134 279648 165218
rect 279328 164898 279370 165134
rect 279606 164898 279648 165134
rect 279328 164866 279648 164898
rect 310048 165454 310368 165486
rect 310048 165218 310090 165454
rect 310326 165218 310368 165454
rect 310048 165134 310368 165218
rect 310048 164898 310090 165134
rect 310326 164898 310368 165134
rect 310048 164866 310368 164898
rect 340768 165454 341088 165486
rect 340768 165218 340810 165454
rect 341046 165218 341088 165454
rect 340768 165134 341088 165218
rect 340768 164898 340810 165134
rect 341046 164898 341088 165134
rect 340768 164866 341088 164898
rect 371488 165454 371808 165486
rect 371488 165218 371530 165454
rect 371766 165218 371808 165454
rect 371488 165134 371808 165218
rect 371488 164898 371530 165134
rect 371766 164898 371808 165134
rect 371488 164866 371808 164898
rect 402208 165454 402528 165486
rect 402208 165218 402250 165454
rect 402486 165218 402528 165454
rect 402208 165134 402528 165218
rect 402208 164898 402250 165134
rect 402486 164898 402528 165134
rect 402208 164866 402528 164898
rect 432928 165454 433248 165486
rect 432928 165218 432970 165454
rect 433206 165218 433248 165454
rect 432928 165134 433248 165218
rect 432928 164898 432970 165134
rect 433206 164898 433248 165134
rect 432928 164866 433248 164898
rect 463648 165454 463968 165486
rect 463648 165218 463690 165454
rect 463926 165218 463968 165454
rect 463648 165134 463968 165218
rect 463648 164898 463690 165134
rect 463926 164898 463968 165134
rect 463648 164866 463968 164898
rect 494368 165454 494688 165486
rect 494368 165218 494410 165454
rect 494646 165218 494688 165454
rect 494368 165134 494688 165218
rect 494368 164898 494410 165134
rect 494646 164898 494688 165134
rect 494368 164866 494688 164898
rect 525088 165454 525408 165486
rect 525088 165218 525130 165454
rect 525366 165218 525408 165454
rect 525088 165134 525408 165218
rect 525088 164898 525130 165134
rect 525366 164898 525408 165134
rect 525088 164866 525408 164898
rect 48928 147454 49248 147486
rect 48928 147218 48970 147454
rect 49206 147218 49248 147454
rect 48928 147134 49248 147218
rect 48928 146898 48970 147134
rect 49206 146898 49248 147134
rect 48928 146866 49248 146898
rect 79648 147454 79968 147486
rect 79648 147218 79690 147454
rect 79926 147218 79968 147454
rect 79648 147134 79968 147218
rect 79648 146898 79690 147134
rect 79926 146898 79968 147134
rect 79648 146866 79968 146898
rect 110368 147454 110688 147486
rect 110368 147218 110410 147454
rect 110646 147218 110688 147454
rect 110368 147134 110688 147218
rect 110368 146898 110410 147134
rect 110646 146898 110688 147134
rect 110368 146866 110688 146898
rect 141088 147454 141408 147486
rect 141088 147218 141130 147454
rect 141366 147218 141408 147454
rect 141088 147134 141408 147218
rect 141088 146898 141130 147134
rect 141366 146898 141408 147134
rect 141088 146866 141408 146898
rect 171808 147454 172128 147486
rect 171808 147218 171850 147454
rect 172086 147218 172128 147454
rect 171808 147134 172128 147218
rect 171808 146898 171850 147134
rect 172086 146898 172128 147134
rect 171808 146866 172128 146898
rect 202528 147454 202848 147486
rect 202528 147218 202570 147454
rect 202806 147218 202848 147454
rect 202528 147134 202848 147218
rect 202528 146898 202570 147134
rect 202806 146898 202848 147134
rect 202528 146866 202848 146898
rect 233248 147454 233568 147486
rect 233248 147218 233290 147454
rect 233526 147218 233568 147454
rect 233248 147134 233568 147218
rect 233248 146898 233290 147134
rect 233526 146898 233568 147134
rect 233248 146866 233568 146898
rect 263968 147454 264288 147486
rect 263968 147218 264010 147454
rect 264246 147218 264288 147454
rect 263968 147134 264288 147218
rect 263968 146898 264010 147134
rect 264246 146898 264288 147134
rect 263968 146866 264288 146898
rect 294688 147454 295008 147486
rect 294688 147218 294730 147454
rect 294966 147218 295008 147454
rect 294688 147134 295008 147218
rect 294688 146898 294730 147134
rect 294966 146898 295008 147134
rect 294688 146866 295008 146898
rect 325408 147454 325728 147486
rect 325408 147218 325450 147454
rect 325686 147218 325728 147454
rect 325408 147134 325728 147218
rect 325408 146898 325450 147134
rect 325686 146898 325728 147134
rect 325408 146866 325728 146898
rect 356128 147454 356448 147486
rect 356128 147218 356170 147454
rect 356406 147218 356448 147454
rect 356128 147134 356448 147218
rect 356128 146898 356170 147134
rect 356406 146898 356448 147134
rect 356128 146866 356448 146898
rect 386848 147454 387168 147486
rect 386848 147218 386890 147454
rect 387126 147218 387168 147454
rect 386848 147134 387168 147218
rect 386848 146898 386890 147134
rect 387126 146898 387168 147134
rect 386848 146866 387168 146898
rect 417568 147454 417888 147486
rect 417568 147218 417610 147454
rect 417846 147218 417888 147454
rect 417568 147134 417888 147218
rect 417568 146898 417610 147134
rect 417846 146898 417888 147134
rect 417568 146866 417888 146898
rect 448288 147454 448608 147486
rect 448288 147218 448330 147454
rect 448566 147218 448608 147454
rect 448288 147134 448608 147218
rect 448288 146898 448330 147134
rect 448566 146898 448608 147134
rect 448288 146866 448608 146898
rect 479008 147454 479328 147486
rect 479008 147218 479050 147454
rect 479286 147218 479328 147454
rect 479008 147134 479328 147218
rect 479008 146898 479050 147134
rect 479286 146898 479328 147134
rect 479008 146866 479328 146898
rect 509728 147454 510048 147486
rect 509728 147218 509770 147454
rect 510006 147218 510048 147454
rect 509728 147134 510048 147218
rect 509728 146898 509770 147134
rect 510006 146898 510048 147134
rect 509728 146866 510048 146898
rect 33568 129454 33888 129486
rect 33568 129218 33610 129454
rect 33846 129218 33888 129454
rect 33568 129134 33888 129218
rect 33568 128898 33610 129134
rect 33846 128898 33888 129134
rect 33568 128866 33888 128898
rect 64288 129454 64608 129486
rect 64288 129218 64330 129454
rect 64566 129218 64608 129454
rect 64288 129134 64608 129218
rect 64288 128898 64330 129134
rect 64566 128898 64608 129134
rect 64288 128866 64608 128898
rect 95008 129454 95328 129486
rect 95008 129218 95050 129454
rect 95286 129218 95328 129454
rect 95008 129134 95328 129218
rect 95008 128898 95050 129134
rect 95286 128898 95328 129134
rect 95008 128866 95328 128898
rect 125728 129454 126048 129486
rect 125728 129218 125770 129454
rect 126006 129218 126048 129454
rect 125728 129134 126048 129218
rect 125728 128898 125770 129134
rect 126006 128898 126048 129134
rect 125728 128866 126048 128898
rect 156448 129454 156768 129486
rect 156448 129218 156490 129454
rect 156726 129218 156768 129454
rect 156448 129134 156768 129218
rect 156448 128898 156490 129134
rect 156726 128898 156768 129134
rect 156448 128866 156768 128898
rect 187168 129454 187488 129486
rect 187168 129218 187210 129454
rect 187446 129218 187488 129454
rect 187168 129134 187488 129218
rect 187168 128898 187210 129134
rect 187446 128898 187488 129134
rect 187168 128866 187488 128898
rect 217888 129454 218208 129486
rect 217888 129218 217930 129454
rect 218166 129218 218208 129454
rect 217888 129134 218208 129218
rect 217888 128898 217930 129134
rect 218166 128898 218208 129134
rect 217888 128866 218208 128898
rect 248608 129454 248928 129486
rect 248608 129218 248650 129454
rect 248886 129218 248928 129454
rect 248608 129134 248928 129218
rect 248608 128898 248650 129134
rect 248886 128898 248928 129134
rect 248608 128866 248928 128898
rect 279328 129454 279648 129486
rect 279328 129218 279370 129454
rect 279606 129218 279648 129454
rect 279328 129134 279648 129218
rect 279328 128898 279370 129134
rect 279606 128898 279648 129134
rect 279328 128866 279648 128898
rect 310048 129454 310368 129486
rect 310048 129218 310090 129454
rect 310326 129218 310368 129454
rect 310048 129134 310368 129218
rect 310048 128898 310090 129134
rect 310326 128898 310368 129134
rect 310048 128866 310368 128898
rect 340768 129454 341088 129486
rect 340768 129218 340810 129454
rect 341046 129218 341088 129454
rect 340768 129134 341088 129218
rect 340768 128898 340810 129134
rect 341046 128898 341088 129134
rect 340768 128866 341088 128898
rect 371488 129454 371808 129486
rect 371488 129218 371530 129454
rect 371766 129218 371808 129454
rect 371488 129134 371808 129218
rect 371488 128898 371530 129134
rect 371766 128898 371808 129134
rect 371488 128866 371808 128898
rect 402208 129454 402528 129486
rect 402208 129218 402250 129454
rect 402486 129218 402528 129454
rect 402208 129134 402528 129218
rect 402208 128898 402250 129134
rect 402486 128898 402528 129134
rect 402208 128866 402528 128898
rect 432928 129454 433248 129486
rect 432928 129218 432970 129454
rect 433206 129218 433248 129454
rect 432928 129134 433248 129218
rect 432928 128898 432970 129134
rect 433206 128898 433248 129134
rect 432928 128866 433248 128898
rect 463648 129454 463968 129486
rect 463648 129218 463690 129454
rect 463926 129218 463968 129454
rect 463648 129134 463968 129218
rect 463648 128898 463690 129134
rect 463926 128898 463968 129134
rect 463648 128866 463968 128898
rect 494368 129454 494688 129486
rect 494368 129218 494410 129454
rect 494646 129218 494688 129454
rect 494368 129134 494688 129218
rect 494368 128898 494410 129134
rect 494646 128898 494688 129134
rect 494368 128866 494688 128898
rect 525088 129454 525408 129486
rect 525088 129218 525130 129454
rect 525366 129218 525408 129454
rect 525088 129134 525408 129218
rect 525088 128898 525130 129134
rect 525366 128898 525408 129134
rect 525088 128866 525408 128898
rect 48928 111454 49248 111486
rect 48928 111218 48970 111454
rect 49206 111218 49248 111454
rect 48928 111134 49248 111218
rect 48928 110898 48970 111134
rect 49206 110898 49248 111134
rect 48928 110866 49248 110898
rect 79648 111454 79968 111486
rect 79648 111218 79690 111454
rect 79926 111218 79968 111454
rect 79648 111134 79968 111218
rect 79648 110898 79690 111134
rect 79926 110898 79968 111134
rect 79648 110866 79968 110898
rect 110368 111454 110688 111486
rect 110368 111218 110410 111454
rect 110646 111218 110688 111454
rect 110368 111134 110688 111218
rect 110368 110898 110410 111134
rect 110646 110898 110688 111134
rect 110368 110866 110688 110898
rect 141088 111454 141408 111486
rect 141088 111218 141130 111454
rect 141366 111218 141408 111454
rect 141088 111134 141408 111218
rect 141088 110898 141130 111134
rect 141366 110898 141408 111134
rect 141088 110866 141408 110898
rect 171808 111454 172128 111486
rect 171808 111218 171850 111454
rect 172086 111218 172128 111454
rect 171808 111134 172128 111218
rect 171808 110898 171850 111134
rect 172086 110898 172128 111134
rect 171808 110866 172128 110898
rect 202528 111454 202848 111486
rect 202528 111218 202570 111454
rect 202806 111218 202848 111454
rect 202528 111134 202848 111218
rect 202528 110898 202570 111134
rect 202806 110898 202848 111134
rect 202528 110866 202848 110898
rect 233248 111454 233568 111486
rect 233248 111218 233290 111454
rect 233526 111218 233568 111454
rect 233248 111134 233568 111218
rect 233248 110898 233290 111134
rect 233526 110898 233568 111134
rect 233248 110866 233568 110898
rect 263968 111454 264288 111486
rect 263968 111218 264010 111454
rect 264246 111218 264288 111454
rect 263968 111134 264288 111218
rect 263968 110898 264010 111134
rect 264246 110898 264288 111134
rect 263968 110866 264288 110898
rect 294688 111454 295008 111486
rect 294688 111218 294730 111454
rect 294966 111218 295008 111454
rect 294688 111134 295008 111218
rect 294688 110898 294730 111134
rect 294966 110898 295008 111134
rect 294688 110866 295008 110898
rect 325408 111454 325728 111486
rect 325408 111218 325450 111454
rect 325686 111218 325728 111454
rect 325408 111134 325728 111218
rect 325408 110898 325450 111134
rect 325686 110898 325728 111134
rect 325408 110866 325728 110898
rect 356128 111454 356448 111486
rect 356128 111218 356170 111454
rect 356406 111218 356448 111454
rect 356128 111134 356448 111218
rect 356128 110898 356170 111134
rect 356406 110898 356448 111134
rect 356128 110866 356448 110898
rect 386848 111454 387168 111486
rect 386848 111218 386890 111454
rect 387126 111218 387168 111454
rect 386848 111134 387168 111218
rect 386848 110898 386890 111134
rect 387126 110898 387168 111134
rect 386848 110866 387168 110898
rect 417568 111454 417888 111486
rect 417568 111218 417610 111454
rect 417846 111218 417888 111454
rect 417568 111134 417888 111218
rect 417568 110898 417610 111134
rect 417846 110898 417888 111134
rect 417568 110866 417888 110898
rect 448288 111454 448608 111486
rect 448288 111218 448330 111454
rect 448566 111218 448608 111454
rect 448288 111134 448608 111218
rect 448288 110898 448330 111134
rect 448566 110898 448608 111134
rect 448288 110866 448608 110898
rect 479008 111454 479328 111486
rect 479008 111218 479050 111454
rect 479286 111218 479328 111454
rect 479008 111134 479328 111218
rect 479008 110898 479050 111134
rect 479286 110898 479328 111134
rect 479008 110866 479328 110898
rect 509728 111454 510048 111486
rect 509728 111218 509770 111454
rect 510006 111218 510048 111454
rect 509728 111134 510048 111218
rect 509728 110898 509770 111134
rect 510006 110898 510048 111134
rect 509728 110866 510048 110898
rect 33568 93454 33888 93486
rect 33568 93218 33610 93454
rect 33846 93218 33888 93454
rect 33568 93134 33888 93218
rect 33568 92898 33610 93134
rect 33846 92898 33888 93134
rect 33568 92866 33888 92898
rect 64288 93454 64608 93486
rect 64288 93218 64330 93454
rect 64566 93218 64608 93454
rect 64288 93134 64608 93218
rect 64288 92898 64330 93134
rect 64566 92898 64608 93134
rect 64288 92866 64608 92898
rect 95008 93454 95328 93486
rect 95008 93218 95050 93454
rect 95286 93218 95328 93454
rect 95008 93134 95328 93218
rect 95008 92898 95050 93134
rect 95286 92898 95328 93134
rect 95008 92866 95328 92898
rect 125728 93454 126048 93486
rect 125728 93218 125770 93454
rect 126006 93218 126048 93454
rect 125728 93134 126048 93218
rect 125728 92898 125770 93134
rect 126006 92898 126048 93134
rect 125728 92866 126048 92898
rect 156448 93454 156768 93486
rect 156448 93218 156490 93454
rect 156726 93218 156768 93454
rect 156448 93134 156768 93218
rect 156448 92898 156490 93134
rect 156726 92898 156768 93134
rect 156448 92866 156768 92898
rect 187168 93454 187488 93486
rect 187168 93218 187210 93454
rect 187446 93218 187488 93454
rect 187168 93134 187488 93218
rect 187168 92898 187210 93134
rect 187446 92898 187488 93134
rect 187168 92866 187488 92898
rect 217888 93454 218208 93486
rect 217888 93218 217930 93454
rect 218166 93218 218208 93454
rect 217888 93134 218208 93218
rect 217888 92898 217930 93134
rect 218166 92898 218208 93134
rect 217888 92866 218208 92898
rect 248608 93454 248928 93486
rect 248608 93218 248650 93454
rect 248886 93218 248928 93454
rect 248608 93134 248928 93218
rect 248608 92898 248650 93134
rect 248886 92898 248928 93134
rect 248608 92866 248928 92898
rect 279328 93454 279648 93486
rect 279328 93218 279370 93454
rect 279606 93218 279648 93454
rect 279328 93134 279648 93218
rect 279328 92898 279370 93134
rect 279606 92898 279648 93134
rect 279328 92866 279648 92898
rect 310048 93454 310368 93486
rect 310048 93218 310090 93454
rect 310326 93218 310368 93454
rect 310048 93134 310368 93218
rect 310048 92898 310090 93134
rect 310326 92898 310368 93134
rect 310048 92866 310368 92898
rect 340768 93454 341088 93486
rect 340768 93218 340810 93454
rect 341046 93218 341088 93454
rect 340768 93134 341088 93218
rect 340768 92898 340810 93134
rect 341046 92898 341088 93134
rect 340768 92866 341088 92898
rect 371488 93454 371808 93486
rect 371488 93218 371530 93454
rect 371766 93218 371808 93454
rect 371488 93134 371808 93218
rect 371488 92898 371530 93134
rect 371766 92898 371808 93134
rect 371488 92866 371808 92898
rect 402208 93454 402528 93486
rect 402208 93218 402250 93454
rect 402486 93218 402528 93454
rect 402208 93134 402528 93218
rect 402208 92898 402250 93134
rect 402486 92898 402528 93134
rect 402208 92866 402528 92898
rect 432928 93454 433248 93486
rect 432928 93218 432970 93454
rect 433206 93218 433248 93454
rect 432928 93134 433248 93218
rect 432928 92898 432970 93134
rect 433206 92898 433248 93134
rect 432928 92866 433248 92898
rect 463648 93454 463968 93486
rect 463648 93218 463690 93454
rect 463926 93218 463968 93454
rect 463648 93134 463968 93218
rect 463648 92898 463690 93134
rect 463926 92898 463968 93134
rect 463648 92866 463968 92898
rect 494368 93454 494688 93486
rect 494368 93218 494410 93454
rect 494646 93218 494688 93454
rect 494368 93134 494688 93218
rect 494368 92898 494410 93134
rect 494646 92898 494688 93134
rect 494368 92866 494688 92898
rect 525088 93454 525408 93486
rect 525088 93218 525130 93454
rect 525366 93218 525408 93454
rect 525088 93134 525408 93218
rect 525088 92898 525130 93134
rect 525366 92898 525408 93134
rect 525088 92866 525408 92898
rect 48928 75454 49248 75486
rect 48928 75218 48970 75454
rect 49206 75218 49248 75454
rect 48928 75134 49248 75218
rect 48928 74898 48970 75134
rect 49206 74898 49248 75134
rect 48928 74866 49248 74898
rect 79648 75454 79968 75486
rect 79648 75218 79690 75454
rect 79926 75218 79968 75454
rect 79648 75134 79968 75218
rect 79648 74898 79690 75134
rect 79926 74898 79968 75134
rect 79648 74866 79968 74898
rect 110368 75454 110688 75486
rect 110368 75218 110410 75454
rect 110646 75218 110688 75454
rect 110368 75134 110688 75218
rect 110368 74898 110410 75134
rect 110646 74898 110688 75134
rect 110368 74866 110688 74898
rect 141088 75454 141408 75486
rect 141088 75218 141130 75454
rect 141366 75218 141408 75454
rect 141088 75134 141408 75218
rect 141088 74898 141130 75134
rect 141366 74898 141408 75134
rect 141088 74866 141408 74898
rect 171808 75454 172128 75486
rect 171808 75218 171850 75454
rect 172086 75218 172128 75454
rect 171808 75134 172128 75218
rect 171808 74898 171850 75134
rect 172086 74898 172128 75134
rect 171808 74866 172128 74898
rect 202528 75454 202848 75486
rect 202528 75218 202570 75454
rect 202806 75218 202848 75454
rect 202528 75134 202848 75218
rect 202528 74898 202570 75134
rect 202806 74898 202848 75134
rect 202528 74866 202848 74898
rect 233248 75454 233568 75486
rect 233248 75218 233290 75454
rect 233526 75218 233568 75454
rect 233248 75134 233568 75218
rect 233248 74898 233290 75134
rect 233526 74898 233568 75134
rect 233248 74866 233568 74898
rect 263968 75454 264288 75486
rect 263968 75218 264010 75454
rect 264246 75218 264288 75454
rect 263968 75134 264288 75218
rect 263968 74898 264010 75134
rect 264246 74898 264288 75134
rect 263968 74866 264288 74898
rect 294688 75454 295008 75486
rect 294688 75218 294730 75454
rect 294966 75218 295008 75454
rect 294688 75134 295008 75218
rect 294688 74898 294730 75134
rect 294966 74898 295008 75134
rect 294688 74866 295008 74898
rect 325408 75454 325728 75486
rect 325408 75218 325450 75454
rect 325686 75218 325728 75454
rect 325408 75134 325728 75218
rect 325408 74898 325450 75134
rect 325686 74898 325728 75134
rect 325408 74866 325728 74898
rect 356128 75454 356448 75486
rect 356128 75218 356170 75454
rect 356406 75218 356448 75454
rect 356128 75134 356448 75218
rect 356128 74898 356170 75134
rect 356406 74898 356448 75134
rect 356128 74866 356448 74898
rect 386848 75454 387168 75486
rect 386848 75218 386890 75454
rect 387126 75218 387168 75454
rect 386848 75134 387168 75218
rect 386848 74898 386890 75134
rect 387126 74898 387168 75134
rect 386848 74866 387168 74898
rect 417568 75454 417888 75486
rect 417568 75218 417610 75454
rect 417846 75218 417888 75454
rect 417568 75134 417888 75218
rect 417568 74898 417610 75134
rect 417846 74898 417888 75134
rect 417568 74866 417888 74898
rect 448288 75454 448608 75486
rect 448288 75218 448330 75454
rect 448566 75218 448608 75454
rect 448288 75134 448608 75218
rect 448288 74898 448330 75134
rect 448566 74898 448608 75134
rect 448288 74866 448608 74898
rect 479008 75454 479328 75486
rect 479008 75218 479050 75454
rect 479286 75218 479328 75454
rect 479008 75134 479328 75218
rect 479008 74898 479050 75134
rect 479286 74898 479328 75134
rect 479008 74866 479328 74898
rect 509728 75454 510048 75486
rect 509728 75218 509770 75454
rect 510006 75218 510048 75454
rect 509728 75134 510048 75218
rect 509728 74898 509770 75134
rect 510006 74898 510048 75134
rect 509728 74866 510048 74898
rect 33568 57454 33888 57486
rect 33568 57218 33610 57454
rect 33846 57218 33888 57454
rect 33568 57134 33888 57218
rect 33568 56898 33610 57134
rect 33846 56898 33888 57134
rect 33568 56866 33888 56898
rect 64288 57454 64608 57486
rect 64288 57218 64330 57454
rect 64566 57218 64608 57454
rect 64288 57134 64608 57218
rect 64288 56898 64330 57134
rect 64566 56898 64608 57134
rect 64288 56866 64608 56898
rect 95008 57454 95328 57486
rect 95008 57218 95050 57454
rect 95286 57218 95328 57454
rect 95008 57134 95328 57218
rect 95008 56898 95050 57134
rect 95286 56898 95328 57134
rect 95008 56866 95328 56898
rect 125728 57454 126048 57486
rect 125728 57218 125770 57454
rect 126006 57218 126048 57454
rect 125728 57134 126048 57218
rect 125728 56898 125770 57134
rect 126006 56898 126048 57134
rect 125728 56866 126048 56898
rect 156448 57454 156768 57486
rect 156448 57218 156490 57454
rect 156726 57218 156768 57454
rect 156448 57134 156768 57218
rect 156448 56898 156490 57134
rect 156726 56898 156768 57134
rect 156448 56866 156768 56898
rect 187168 57454 187488 57486
rect 187168 57218 187210 57454
rect 187446 57218 187488 57454
rect 187168 57134 187488 57218
rect 187168 56898 187210 57134
rect 187446 56898 187488 57134
rect 187168 56866 187488 56898
rect 217888 57454 218208 57486
rect 217888 57218 217930 57454
rect 218166 57218 218208 57454
rect 217888 57134 218208 57218
rect 217888 56898 217930 57134
rect 218166 56898 218208 57134
rect 217888 56866 218208 56898
rect 248608 57454 248928 57486
rect 248608 57218 248650 57454
rect 248886 57218 248928 57454
rect 248608 57134 248928 57218
rect 248608 56898 248650 57134
rect 248886 56898 248928 57134
rect 248608 56866 248928 56898
rect 279328 57454 279648 57486
rect 279328 57218 279370 57454
rect 279606 57218 279648 57454
rect 279328 57134 279648 57218
rect 279328 56898 279370 57134
rect 279606 56898 279648 57134
rect 279328 56866 279648 56898
rect 310048 57454 310368 57486
rect 310048 57218 310090 57454
rect 310326 57218 310368 57454
rect 310048 57134 310368 57218
rect 310048 56898 310090 57134
rect 310326 56898 310368 57134
rect 310048 56866 310368 56898
rect 340768 57454 341088 57486
rect 340768 57218 340810 57454
rect 341046 57218 341088 57454
rect 340768 57134 341088 57218
rect 340768 56898 340810 57134
rect 341046 56898 341088 57134
rect 340768 56866 341088 56898
rect 371488 57454 371808 57486
rect 371488 57218 371530 57454
rect 371766 57218 371808 57454
rect 371488 57134 371808 57218
rect 371488 56898 371530 57134
rect 371766 56898 371808 57134
rect 371488 56866 371808 56898
rect 402208 57454 402528 57486
rect 402208 57218 402250 57454
rect 402486 57218 402528 57454
rect 402208 57134 402528 57218
rect 402208 56898 402250 57134
rect 402486 56898 402528 57134
rect 402208 56866 402528 56898
rect 432928 57454 433248 57486
rect 432928 57218 432970 57454
rect 433206 57218 433248 57454
rect 432928 57134 433248 57218
rect 432928 56898 432970 57134
rect 433206 56898 433248 57134
rect 432928 56866 433248 56898
rect 463648 57454 463968 57486
rect 463648 57218 463690 57454
rect 463926 57218 463968 57454
rect 463648 57134 463968 57218
rect 463648 56898 463690 57134
rect 463926 56898 463968 57134
rect 463648 56866 463968 56898
rect 494368 57454 494688 57486
rect 494368 57218 494410 57454
rect 494646 57218 494688 57454
rect 494368 57134 494688 57218
rect 494368 56898 494410 57134
rect 494646 56898 494688 57134
rect 494368 56866 494688 56898
rect 525088 57454 525408 57486
rect 525088 57218 525130 57454
rect 525366 57218 525408 57454
rect 525088 57134 525408 57218
rect 525088 56898 525130 57134
rect 525366 56898 525408 57134
rect 525088 56866 525408 56898
rect 30787 45660 30853 45661
rect 30787 45596 30788 45660
rect 30852 45596 30853 45660
rect 30787 45595 30853 45596
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 26003 19412 26069 19413
rect 26003 19348 26004 19412
rect 26068 19348 26069 19412
rect 26003 19347 26069 19348
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 32614 31574 48000
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 39454 38414 48000
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 43174 42134 48000
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 46894 45854 48000
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 48000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 48000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 48000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 48000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 48000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 48000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 48000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 48000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 48000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 48000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 48000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 48000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 48000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 48000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 48000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 48000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 48000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 48000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 48000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 48000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 48000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 48000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 48000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 48000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 48000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 48000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 48000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 48000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 48000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 48000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 48000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 48000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 48000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 48000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 48000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 48000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 48000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 48000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 48000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 48000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 48000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 48000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 48000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 48000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 48000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 48000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 48000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 48000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 48000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 48000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 48000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 48000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 48000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 48000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 48000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 48000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 48000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 48000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 48000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 48000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 48000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 48000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 48000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 48000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 48000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 48000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 48000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 48000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 48000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 48000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 43174 366134 48000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 48000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 48000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 48000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 48000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 48000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 48000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 48000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 48000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 48000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 48000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 48000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 48000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 48000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 48000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 48000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 48000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 48000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 48000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 48000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 48000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 48000
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 48000
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 48000
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 48000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 48000
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 48000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 48000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 48000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 48000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 48000
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 48000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 48000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 48000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 48000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 48000
rect 527222 44301 527282 669291
rect 527219 44300 527285 44301
rect 527219 44236 527220 44300
rect 527284 44236 527285 44300
rect 527219 44235 527285 44236
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 48000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 28894 531854 48000
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 32614 535574 48000
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 536790 31925 536850 669291
rect 540099 667996 540165 667997
rect 540099 667932 540100 667996
rect 540164 667932 540165 667996
rect 540099 667931 540165 667932
rect 540102 484618 540162 667931
rect 540448 651454 540768 651486
rect 540448 651218 540490 651454
rect 540726 651218 540768 651454
rect 540448 651134 540768 651218
rect 540448 650898 540490 651134
rect 540726 650898 540768 651134
rect 540448 650866 540768 650898
rect 540448 615454 540768 615486
rect 540448 615218 540490 615454
rect 540726 615218 540768 615454
rect 540448 615134 540768 615218
rect 540448 614898 540490 615134
rect 540726 614898 540768 615134
rect 540448 614866 540768 614898
rect 540448 579454 540768 579486
rect 540448 579218 540490 579454
rect 540726 579218 540768 579454
rect 540448 579134 540768 579218
rect 540448 578898 540490 579134
rect 540726 578898 540768 579134
rect 540448 578866 540768 578898
rect 540448 543454 540768 543486
rect 540448 543218 540490 543454
rect 540726 543218 540768 543454
rect 540448 543134 540768 543218
rect 540448 542898 540490 543134
rect 540726 542898 540768 543134
rect 540448 542866 540768 542898
rect 540448 507454 540768 507486
rect 540448 507218 540490 507454
rect 540726 507218 540768 507454
rect 540448 507134 540768 507218
rect 540448 506898 540490 507134
rect 540726 506898 540768 507134
rect 540448 506866 540768 506898
rect 541022 499590 541082 669291
rect 541022 499530 541450 499590
rect 540448 471454 540768 471486
rect 540448 471218 540490 471454
rect 540726 471218 540768 471454
rect 540448 471134 540768 471218
rect 540448 470898 540490 471134
rect 540726 470898 540768 471134
rect 540448 470866 540768 470898
rect 541390 470610 541450 499530
rect 541022 470550 541450 470610
rect 540448 435454 540768 435486
rect 540448 435218 540490 435454
rect 540726 435218 540768 435454
rect 540448 435134 540768 435218
rect 540448 434898 540490 435134
rect 540726 434898 540768 435134
rect 540448 434866 540768 434898
rect 540448 399454 540768 399486
rect 540448 399218 540490 399454
rect 540726 399218 540768 399454
rect 540448 399134 540768 399218
rect 540448 398898 540490 399134
rect 540726 398898 540768 399134
rect 540448 398866 540768 398898
rect 540448 363454 540768 363486
rect 540448 363218 540490 363454
rect 540726 363218 540768 363454
rect 540448 363134 540768 363218
rect 540448 362898 540490 363134
rect 540726 362898 540768 363134
rect 540448 362866 540768 362898
rect 540448 327454 540768 327486
rect 540448 327218 540490 327454
rect 540726 327218 540768 327454
rect 540448 327134 540768 327218
rect 540448 326898 540490 327134
rect 540726 326898 540768 327134
rect 540448 326866 540768 326898
rect 540448 291454 540768 291486
rect 540448 291218 540490 291454
rect 540726 291218 540768 291454
rect 540448 291134 540768 291218
rect 540448 290898 540490 291134
rect 540726 290898 540768 291134
rect 540448 290866 540768 290898
rect 540448 255454 540768 255486
rect 540448 255218 540490 255454
rect 540726 255218 540768 255454
rect 540448 255134 540768 255218
rect 540448 254898 540490 255134
rect 540726 254898 540768 255134
rect 540448 254866 540768 254898
rect 540448 219454 540768 219486
rect 540448 219218 540490 219454
rect 540726 219218 540768 219454
rect 540448 219134 540768 219218
rect 540448 218898 540490 219134
rect 540726 218898 540768 219134
rect 540448 218866 540768 218898
rect 540448 183454 540768 183486
rect 540448 183218 540490 183454
rect 540726 183218 540768 183454
rect 540448 183134 540768 183218
rect 540448 182898 540490 183134
rect 540726 182898 540768 183134
rect 540448 182866 540768 182898
rect 540448 147454 540768 147486
rect 540448 147218 540490 147454
rect 540726 147218 540768 147454
rect 540448 147134 540768 147218
rect 540448 146898 540490 147134
rect 540726 146898 540768 147134
rect 540448 146866 540768 146898
rect 540448 111454 540768 111486
rect 540448 111218 540490 111454
rect 540726 111218 540768 111454
rect 540448 111134 540768 111218
rect 540448 110898 540490 111134
rect 540726 110898 540768 111134
rect 540448 110866 540768 110898
rect 540448 75454 540768 75486
rect 540448 75218 540490 75454
rect 540726 75218 540768 75454
rect 540448 75134 540768 75218
rect 540448 74898 540490 75134
rect 540726 74898 540768 75134
rect 540448 74866 540768 74898
rect 536787 31924 536853 31925
rect 536787 31860 536788 31924
rect 536852 31860 536853 31924
rect 536787 31859 536853 31860
rect 541022 5813 541082 470550
rect 541794 39454 542414 48000
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541019 5812 541085 5813
rect 541019 5748 541020 5812
rect 541084 5748 541085 5812
rect 541019 5747 541085 5748
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 43174 546134 48000
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 546542 19549 546602 669291
rect 553902 71909 553962 669427
rect 554086 85645 554146 670787
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 554083 85644 554149 85645
rect 554083 85580 554084 85644
rect 554148 85580 554149 85644
rect 554083 85579 554149 85580
rect 553899 71908 553965 71909
rect 553899 71844 553900 71908
rect 553964 71844 553965 71908
rect 553899 71843 553965 71844
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 549234 46894 549854 48000
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 546539 19548 546605 19549
rect 546539 19484 546540 19548
rect 546604 19484 546605 19548
rect 546539 19483 546605 19484
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 14614 553574 48000
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 18250 651218 18486 651454
rect 18250 650898 18486 651134
rect 18250 615218 18486 615454
rect 18250 614898 18486 615134
rect 18250 579218 18486 579454
rect 18250 578898 18486 579134
rect 18250 543218 18486 543454
rect 18250 542898 18486 543134
rect 18250 507218 18486 507454
rect 18250 506898 18486 507134
rect 18250 471218 18486 471454
rect 18250 470898 18486 471134
rect 18250 435218 18486 435454
rect 18250 434898 18486 435134
rect 18250 399218 18486 399454
rect 18250 398898 18486 399134
rect 18250 363218 18486 363454
rect 18250 362898 18486 363134
rect 18250 327218 18486 327454
rect 18250 326898 18486 327134
rect 18250 291218 18486 291454
rect 18250 290898 18486 291134
rect 18250 255218 18486 255454
rect 18250 254898 18486 255134
rect 18250 219218 18486 219454
rect 18250 218898 18486 219134
rect 18250 183218 18486 183454
rect 18250 182898 18486 183134
rect 18250 147218 18486 147454
rect 18250 146898 18486 147134
rect 18250 111218 18486 111454
rect 18250 110898 18486 111134
rect 18250 75218 18486 75454
rect 18250 74898 18486 75134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 48970 651218 49206 651454
rect 48970 650898 49206 651134
rect 79690 651218 79926 651454
rect 79690 650898 79926 651134
rect 110410 651218 110646 651454
rect 110410 650898 110646 651134
rect 141130 651218 141366 651454
rect 141130 650898 141366 651134
rect 171850 651218 172086 651454
rect 171850 650898 172086 651134
rect 202570 651218 202806 651454
rect 202570 650898 202806 651134
rect 233290 651218 233526 651454
rect 233290 650898 233526 651134
rect 264010 651218 264246 651454
rect 264010 650898 264246 651134
rect 294730 651218 294966 651454
rect 294730 650898 294966 651134
rect 325450 651218 325686 651454
rect 325450 650898 325686 651134
rect 356170 651218 356406 651454
rect 356170 650898 356406 651134
rect 386890 651218 387126 651454
rect 386890 650898 387126 651134
rect 417610 651218 417846 651454
rect 417610 650898 417846 651134
rect 448330 651218 448566 651454
rect 448330 650898 448566 651134
rect 479050 651218 479286 651454
rect 479050 650898 479286 651134
rect 509770 651218 510006 651454
rect 509770 650898 510006 651134
rect 33610 633218 33846 633454
rect 33610 632898 33846 633134
rect 64330 633218 64566 633454
rect 64330 632898 64566 633134
rect 95050 633218 95286 633454
rect 95050 632898 95286 633134
rect 125770 633218 126006 633454
rect 125770 632898 126006 633134
rect 156490 633218 156726 633454
rect 156490 632898 156726 633134
rect 187210 633218 187446 633454
rect 187210 632898 187446 633134
rect 217930 633218 218166 633454
rect 217930 632898 218166 633134
rect 248650 633218 248886 633454
rect 248650 632898 248886 633134
rect 279370 633218 279606 633454
rect 279370 632898 279606 633134
rect 310090 633218 310326 633454
rect 310090 632898 310326 633134
rect 340810 633218 341046 633454
rect 340810 632898 341046 633134
rect 371530 633218 371766 633454
rect 371530 632898 371766 633134
rect 402250 633218 402486 633454
rect 402250 632898 402486 633134
rect 432970 633218 433206 633454
rect 432970 632898 433206 633134
rect 463690 633218 463926 633454
rect 463690 632898 463926 633134
rect 494410 633218 494646 633454
rect 494410 632898 494646 633134
rect 525130 633218 525366 633454
rect 525130 632898 525366 633134
rect 48970 615218 49206 615454
rect 48970 614898 49206 615134
rect 79690 615218 79926 615454
rect 79690 614898 79926 615134
rect 110410 615218 110646 615454
rect 110410 614898 110646 615134
rect 141130 615218 141366 615454
rect 141130 614898 141366 615134
rect 171850 615218 172086 615454
rect 171850 614898 172086 615134
rect 202570 615218 202806 615454
rect 202570 614898 202806 615134
rect 233290 615218 233526 615454
rect 233290 614898 233526 615134
rect 264010 615218 264246 615454
rect 264010 614898 264246 615134
rect 294730 615218 294966 615454
rect 294730 614898 294966 615134
rect 325450 615218 325686 615454
rect 325450 614898 325686 615134
rect 356170 615218 356406 615454
rect 356170 614898 356406 615134
rect 386890 615218 387126 615454
rect 386890 614898 387126 615134
rect 417610 615218 417846 615454
rect 417610 614898 417846 615134
rect 448330 615218 448566 615454
rect 448330 614898 448566 615134
rect 479050 615218 479286 615454
rect 479050 614898 479286 615134
rect 509770 615218 510006 615454
rect 509770 614898 510006 615134
rect 33610 597218 33846 597454
rect 33610 596898 33846 597134
rect 64330 597218 64566 597454
rect 64330 596898 64566 597134
rect 95050 597218 95286 597454
rect 95050 596898 95286 597134
rect 125770 597218 126006 597454
rect 125770 596898 126006 597134
rect 156490 597218 156726 597454
rect 156490 596898 156726 597134
rect 187210 597218 187446 597454
rect 187210 596898 187446 597134
rect 217930 597218 218166 597454
rect 217930 596898 218166 597134
rect 248650 597218 248886 597454
rect 248650 596898 248886 597134
rect 279370 597218 279606 597454
rect 279370 596898 279606 597134
rect 310090 597218 310326 597454
rect 310090 596898 310326 597134
rect 340810 597218 341046 597454
rect 340810 596898 341046 597134
rect 371530 597218 371766 597454
rect 371530 596898 371766 597134
rect 402250 597218 402486 597454
rect 402250 596898 402486 597134
rect 432970 597218 433206 597454
rect 432970 596898 433206 597134
rect 463690 597218 463926 597454
rect 463690 596898 463926 597134
rect 494410 597218 494646 597454
rect 494410 596898 494646 597134
rect 525130 597218 525366 597454
rect 525130 596898 525366 597134
rect 48970 579218 49206 579454
rect 48970 578898 49206 579134
rect 79690 579218 79926 579454
rect 79690 578898 79926 579134
rect 110410 579218 110646 579454
rect 110410 578898 110646 579134
rect 141130 579218 141366 579454
rect 141130 578898 141366 579134
rect 171850 579218 172086 579454
rect 171850 578898 172086 579134
rect 202570 579218 202806 579454
rect 202570 578898 202806 579134
rect 233290 579218 233526 579454
rect 233290 578898 233526 579134
rect 264010 579218 264246 579454
rect 264010 578898 264246 579134
rect 294730 579218 294966 579454
rect 294730 578898 294966 579134
rect 325450 579218 325686 579454
rect 325450 578898 325686 579134
rect 356170 579218 356406 579454
rect 356170 578898 356406 579134
rect 386890 579218 387126 579454
rect 386890 578898 387126 579134
rect 417610 579218 417846 579454
rect 417610 578898 417846 579134
rect 448330 579218 448566 579454
rect 448330 578898 448566 579134
rect 479050 579218 479286 579454
rect 479050 578898 479286 579134
rect 509770 579218 510006 579454
rect 509770 578898 510006 579134
rect 33610 561218 33846 561454
rect 33610 560898 33846 561134
rect 64330 561218 64566 561454
rect 64330 560898 64566 561134
rect 95050 561218 95286 561454
rect 95050 560898 95286 561134
rect 125770 561218 126006 561454
rect 125770 560898 126006 561134
rect 156490 561218 156726 561454
rect 156490 560898 156726 561134
rect 187210 561218 187446 561454
rect 187210 560898 187446 561134
rect 217930 561218 218166 561454
rect 217930 560898 218166 561134
rect 248650 561218 248886 561454
rect 248650 560898 248886 561134
rect 279370 561218 279606 561454
rect 279370 560898 279606 561134
rect 310090 561218 310326 561454
rect 310090 560898 310326 561134
rect 340810 561218 341046 561454
rect 340810 560898 341046 561134
rect 371530 561218 371766 561454
rect 371530 560898 371766 561134
rect 402250 561218 402486 561454
rect 402250 560898 402486 561134
rect 432970 561218 433206 561454
rect 432970 560898 433206 561134
rect 463690 561218 463926 561454
rect 463690 560898 463926 561134
rect 494410 561218 494646 561454
rect 494410 560898 494646 561134
rect 525130 561218 525366 561454
rect 525130 560898 525366 561134
rect 48970 543218 49206 543454
rect 48970 542898 49206 543134
rect 79690 543218 79926 543454
rect 79690 542898 79926 543134
rect 110410 543218 110646 543454
rect 110410 542898 110646 543134
rect 141130 543218 141366 543454
rect 141130 542898 141366 543134
rect 171850 543218 172086 543454
rect 171850 542898 172086 543134
rect 202570 543218 202806 543454
rect 202570 542898 202806 543134
rect 233290 543218 233526 543454
rect 233290 542898 233526 543134
rect 264010 543218 264246 543454
rect 264010 542898 264246 543134
rect 294730 543218 294966 543454
rect 294730 542898 294966 543134
rect 325450 543218 325686 543454
rect 325450 542898 325686 543134
rect 356170 543218 356406 543454
rect 356170 542898 356406 543134
rect 386890 543218 387126 543454
rect 386890 542898 387126 543134
rect 417610 543218 417846 543454
rect 417610 542898 417846 543134
rect 448330 543218 448566 543454
rect 448330 542898 448566 543134
rect 479050 543218 479286 543454
rect 479050 542898 479286 543134
rect 509770 543218 510006 543454
rect 509770 542898 510006 543134
rect 33610 525218 33846 525454
rect 33610 524898 33846 525134
rect 64330 525218 64566 525454
rect 64330 524898 64566 525134
rect 95050 525218 95286 525454
rect 95050 524898 95286 525134
rect 125770 525218 126006 525454
rect 125770 524898 126006 525134
rect 156490 525218 156726 525454
rect 156490 524898 156726 525134
rect 187210 525218 187446 525454
rect 187210 524898 187446 525134
rect 217930 525218 218166 525454
rect 217930 524898 218166 525134
rect 248650 525218 248886 525454
rect 248650 524898 248886 525134
rect 279370 525218 279606 525454
rect 279370 524898 279606 525134
rect 310090 525218 310326 525454
rect 310090 524898 310326 525134
rect 340810 525218 341046 525454
rect 340810 524898 341046 525134
rect 371530 525218 371766 525454
rect 371530 524898 371766 525134
rect 402250 525218 402486 525454
rect 402250 524898 402486 525134
rect 432970 525218 433206 525454
rect 432970 524898 433206 525134
rect 463690 525218 463926 525454
rect 463690 524898 463926 525134
rect 494410 525218 494646 525454
rect 494410 524898 494646 525134
rect 525130 525218 525366 525454
rect 525130 524898 525366 525134
rect 48970 507218 49206 507454
rect 48970 506898 49206 507134
rect 79690 507218 79926 507454
rect 79690 506898 79926 507134
rect 110410 507218 110646 507454
rect 110410 506898 110646 507134
rect 141130 507218 141366 507454
rect 141130 506898 141366 507134
rect 171850 507218 172086 507454
rect 171850 506898 172086 507134
rect 202570 507218 202806 507454
rect 202570 506898 202806 507134
rect 233290 507218 233526 507454
rect 233290 506898 233526 507134
rect 264010 507218 264246 507454
rect 264010 506898 264246 507134
rect 294730 507218 294966 507454
rect 294730 506898 294966 507134
rect 325450 507218 325686 507454
rect 325450 506898 325686 507134
rect 356170 507218 356406 507454
rect 356170 506898 356406 507134
rect 386890 507218 387126 507454
rect 386890 506898 387126 507134
rect 417610 507218 417846 507454
rect 417610 506898 417846 507134
rect 448330 507218 448566 507454
rect 448330 506898 448566 507134
rect 479050 507218 479286 507454
rect 479050 506898 479286 507134
rect 509770 507218 510006 507454
rect 509770 506898 510006 507134
rect 33610 489218 33846 489454
rect 33610 488898 33846 489134
rect 64330 489218 64566 489454
rect 64330 488898 64566 489134
rect 95050 489218 95286 489454
rect 95050 488898 95286 489134
rect 125770 489218 126006 489454
rect 125770 488898 126006 489134
rect 156490 489218 156726 489454
rect 156490 488898 156726 489134
rect 187210 489218 187446 489454
rect 187210 488898 187446 489134
rect 217930 489218 218166 489454
rect 217930 488898 218166 489134
rect 248650 489218 248886 489454
rect 248650 488898 248886 489134
rect 279370 489218 279606 489454
rect 279370 488898 279606 489134
rect 310090 489218 310326 489454
rect 310090 488898 310326 489134
rect 340810 489218 341046 489454
rect 340810 488898 341046 489134
rect 371530 489218 371766 489454
rect 371530 488898 371766 489134
rect 402250 489218 402486 489454
rect 402250 488898 402486 489134
rect 432970 489218 433206 489454
rect 432970 488898 433206 489134
rect 463690 489218 463926 489454
rect 463690 488898 463926 489134
rect 494410 489218 494646 489454
rect 494410 488898 494646 489134
rect 525130 489218 525366 489454
rect 525130 488898 525366 489134
rect 48970 471218 49206 471454
rect 48970 470898 49206 471134
rect 79690 471218 79926 471454
rect 79690 470898 79926 471134
rect 110410 471218 110646 471454
rect 110410 470898 110646 471134
rect 141130 471218 141366 471454
rect 141130 470898 141366 471134
rect 171850 471218 172086 471454
rect 171850 470898 172086 471134
rect 202570 471218 202806 471454
rect 202570 470898 202806 471134
rect 233290 471218 233526 471454
rect 233290 470898 233526 471134
rect 264010 471218 264246 471454
rect 264010 470898 264246 471134
rect 294730 471218 294966 471454
rect 294730 470898 294966 471134
rect 325450 471218 325686 471454
rect 325450 470898 325686 471134
rect 356170 471218 356406 471454
rect 356170 470898 356406 471134
rect 386890 471218 387126 471454
rect 386890 470898 387126 471134
rect 417610 471218 417846 471454
rect 417610 470898 417846 471134
rect 448330 471218 448566 471454
rect 448330 470898 448566 471134
rect 479050 471218 479286 471454
rect 479050 470898 479286 471134
rect 509770 471218 510006 471454
rect 509770 470898 510006 471134
rect 33610 453218 33846 453454
rect 33610 452898 33846 453134
rect 64330 453218 64566 453454
rect 64330 452898 64566 453134
rect 95050 453218 95286 453454
rect 95050 452898 95286 453134
rect 125770 453218 126006 453454
rect 125770 452898 126006 453134
rect 156490 453218 156726 453454
rect 156490 452898 156726 453134
rect 187210 453218 187446 453454
rect 187210 452898 187446 453134
rect 217930 453218 218166 453454
rect 217930 452898 218166 453134
rect 248650 453218 248886 453454
rect 248650 452898 248886 453134
rect 279370 453218 279606 453454
rect 279370 452898 279606 453134
rect 310090 453218 310326 453454
rect 310090 452898 310326 453134
rect 340810 453218 341046 453454
rect 340810 452898 341046 453134
rect 371530 453218 371766 453454
rect 371530 452898 371766 453134
rect 402250 453218 402486 453454
rect 402250 452898 402486 453134
rect 432970 453218 433206 453454
rect 432970 452898 433206 453134
rect 463690 453218 463926 453454
rect 463690 452898 463926 453134
rect 494410 453218 494646 453454
rect 494410 452898 494646 453134
rect 525130 453218 525366 453454
rect 525130 452898 525366 453134
rect 48970 435218 49206 435454
rect 48970 434898 49206 435134
rect 79690 435218 79926 435454
rect 79690 434898 79926 435134
rect 110410 435218 110646 435454
rect 110410 434898 110646 435134
rect 141130 435218 141366 435454
rect 141130 434898 141366 435134
rect 171850 435218 172086 435454
rect 171850 434898 172086 435134
rect 202570 435218 202806 435454
rect 202570 434898 202806 435134
rect 233290 435218 233526 435454
rect 233290 434898 233526 435134
rect 264010 435218 264246 435454
rect 264010 434898 264246 435134
rect 294730 435218 294966 435454
rect 294730 434898 294966 435134
rect 325450 435218 325686 435454
rect 325450 434898 325686 435134
rect 356170 435218 356406 435454
rect 356170 434898 356406 435134
rect 386890 435218 387126 435454
rect 386890 434898 387126 435134
rect 417610 435218 417846 435454
rect 417610 434898 417846 435134
rect 448330 435218 448566 435454
rect 448330 434898 448566 435134
rect 479050 435218 479286 435454
rect 479050 434898 479286 435134
rect 509770 435218 510006 435454
rect 509770 434898 510006 435134
rect 33610 417218 33846 417454
rect 33610 416898 33846 417134
rect 64330 417218 64566 417454
rect 64330 416898 64566 417134
rect 95050 417218 95286 417454
rect 95050 416898 95286 417134
rect 125770 417218 126006 417454
rect 125770 416898 126006 417134
rect 156490 417218 156726 417454
rect 156490 416898 156726 417134
rect 187210 417218 187446 417454
rect 187210 416898 187446 417134
rect 217930 417218 218166 417454
rect 217930 416898 218166 417134
rect 248650 417218 248886 417454
rect 248650 416898 248886 417134
rect 279370 417218 279606 417454
rect 279370 416898 279606 417134
rect 310090 417218 310326 417454
rect 310090 416898 310326 417134
rect 340810 417218 341046 417454
rect 340810 416898 341046 417134
rect 371530 417218 371766 417454
rect 371530 416898 371766 417134
rect 402250 417218 402486 417454
rect 402250 416898 402486 417134
rect 432970 417218 433206 417454
rect 432970 416898 433206 417134
rect 463690 417218 463926 417454
rect 463690 416898 463926 417134
rect 494410 417218 494646 417454
rect 494410 416898 494646 417134
rect 525130 417218 525366 417454
rect 525130 416898 525366 417134
rect 48970 399218 49206 399454
rect 48970 398898 49206 399134
rect 79690 399218 79926 399454
rect 79690 398898 79926 399134
rect 110410 399218 110646 399454
rect 110410 398898 110646 399134
rect 141130 399218 141366 399454
rect 141130 398898 141366 399134
rect 171850 399218 172086 399454
rect 171850 398898 172086 399134
rect 202570 399218 202806 399454
rect 202570 398898 202806 399134
rect 233290 399218 233526 399454
rect 233290 398898 233526 399134
rect 264010 399218 264246 399454
rect 264010 398898 264246 399134
rect 294730 399218 294966 399454
rect 294730 398898 294966 399134
rect 325450 399218 325686 399454
rect 325450 398898 325686 399134
rect 356170 399218 356406 399454
rect 356170 398898 356406 399134
rect 386890 399218 387126 399454
rect 386890 398898 387126 399134
rect 417610 399218 417846 399454
rect 417610 398898 417846 399134
rect 448330 399218 448566 399454
rect 448330 398898 448566 399134
rect 479050 399218 479286 399454
rect 479050 398898 479286 399134
rect 509770 399218 510006 399454
rect 509770 398898 510006 399134
rect 33610 381218 33846 381454
rect 33610 380898 33846 381134
rect 64330 381218 64566 381454
rect 64330 380898 64566 381134
rect 95050 381218 95286 381454
rect 95050 380898 95286 381134
rect 125770 381218 126006 381454
rect 125770 380898 126006 381134
rect 156490 381218 156726 381454
rect 156490 380898 156726 381134
rect 187210 381218 187446 381454
rect 187210 380898 187446 381134
rect 217930 381218 218166 381454
rect 217930 380898 218166 381134
rect 248650 381218 248886 381454
rect 248650 380898 248886 381134
rect 279370 381218 279606 381454
rect 279370 380898 279606 381134
rect 310090 381218 310326 381454
rect 310090 380898 310326 381134
rect 340810 381218 341046 381454
rect 340810 380898 341046 381134
rect 371530 381218 371766 381454
rect 371530 380898 371766 381134
rect 402250 381218 402486 381454
rect 402250 380898 402486 381134
rect 432970 381218 433206 381454
rect 432970 380898 433206 381134
rect 463690 381218 463926 381454
rect 463690 380898 463926 381134
rect 494410 381218 494646 381454
rect 494410 380898 494646 381134
rect 525130 381218 525366 381454
rect 525130 380898 525366 381134
rect 48970 363218 49206 363454
rect 48970 362898 49206 363134
rect 79690 363218 79926 363454
rect 79690 362898 79926 363134
rect 110410 363218 110646 363454
rect 110410 362898 110646 363134
rect 141130 363218 141366 363454
rect 141130 362898 141366 363134
rect 171850 363218 172086 363454
rect 171850 362898 172086 363134
rect 202570 363218 202806 363454
rect 202570 362898 202806 363134
rect 233290 363218 233526 363454
rect 233290 362898 233526 363134
rect 264010 363218 264246 363454
rect 264010 362898 264246 363134
rect 294730 363218 294966 363454
rect 294730 362898 294966 363134
rect 325450 363218 325686 363454
rect 325450 362898 325686 363134
rect 356170 363218 356406 363454
rect 356170 362898 356406 363134
rect 386890 363218 387126 363454
rect 386890 362898 387126 363134
rect 417610 363218 417846 363454
rect 417610 362898 417846 363134
rect 448330 363218 448566 363454
rect 448330 362898 448566 363134
rect 479050 363218 479286 363454
rect 479050 362898 479286 363134
rect 509770 363218 510006 363454
rect 509770 362898 510006 363134
rect 33610 345218 33846 345454
rect 33610 344898 33846 345134
rect 64330 345218 64566 345454
rect 64330 344898 64566 345134
rect 95050 345218 95286 345454
rect 95050 344898 95286 345134
rect 125770 345218 126006 345454
rect 125770 344898 126006 345134
rect 156490 345218 156726 345454
rect 156490 344898 156726 345134
rect 187210 345218 187446 345454
rect 187210 344898 187446 345134
rect 217930 345218 218166 345454
rect 217930 344898 218166 345134
rect 248650 345218 248886 345454
rect 248650 344898 248886 345134
rect 279370 345218 279606 345454
rect 279370 344898 279606 345134
rect 310090 345218 310326 345454
rect 310090 344898 310326 345134
rect 340810 345218 341046 345454
rect 340810 344898 341046 345134
rect 371530 345218 371766 345454
rect 371530 344898 371766 345134
rect 402250 345218 402486 345454
rect 402250 344898 402486 345134
rect 432970 345218 433206 345454
rect 432970 344898 433206 345134
rect 463690 345218 463926 345454
rect 463690 344898 463926 345134
rect 494410 345218 494646 345454
rect 494410 344898 494646 345134
rect 525130 345218 525366 345454
rect 525130 344898 525366 345134
rect 48970 327218 49206 327454
rect 48970 326898 49206 327134
rect 79690 327218 79926 327454
rect 79690 326898 79926 327134
rect 110410 327218 110646 327454
rect 110410 326898 110646 327134
rect 141130 327218 141366 327454
rect 141130 326898 141366 327134
rect 171850 327218 172086 327454
rect 171850 326898 172086 327134
rect 202570 327218 202806 327454
rect 202570 326898 202806 327134
rect 233290 327218 233526 327454
rect 233290 326898 233526 327134
rect 264010 327218 264246 327454
rect 264010 326898 264246 327134
rect 294730 327218 294966 327454
rect 294730 326898 294966 327134
rect 325450 327218 325686 327454
rect 325450 326898 325686 327134
rect 356170 327218 356406 327454
rect 356170 326898 356406 327134
rect 386890 327218 387126 327454
rect 386890 326898 387126 327134
rect 417610 327218 417846 327454
rect 417610 326898 417846 327134
rect 448330 327218 448566 327454
rect 448330 326898 448566 327134
rect 479050 327218 479286 327454
rect 479050 326898 479286 327134
rect 509770 327218 510006 327454
rect 509770 326898 510006 327134
rect 33610 309218 33846 309454
rect 33610 308898 33846 309134
rect 64330 309218 64566 309454
rect 64330 308898 64566 309134
rect 95050 309218 95286 309454
rect 95050 308898 95286 309134
rect 125770 309218 126006 309454
rect 125770 308898 126006 309134
rect 156490 309218 156726 309454
rect 156490 308898 156726 309134
rect 187210 309218 187446 309454
rect 187210 308898 187446 309134
rect 217930 309218 218166 309454
rect 217930 308898 218166 309134
rect 248650 309218 248886 309454
rect 248650 308898 248886 309134
rect 279370 309218 279606 309454
rect 279370 308898 279606 309134
rect 310090 309218 310326 309454
rect 310090 308898 310326 309134
rect 340810 309218 341046 309454
rect 340810 308898 341046 309134
rect 371530 309218 371766 309454
rect 371530 308898 371766 309134
rect 402250 309218 402486 309454
rect 402250 308898 402486 309134
rect 432970 309218 433206 309454
rect 432970 308898 433206 309134
rect 463690 309218 463926 309454
rect 463690 308898 463926 309134
rect 494410 309218 494646 309454
rect 494410 308898 494646 309134
rect 525130 309218 525366 309454
rect 525130 308898 525366 309134
rect 48970 291218 49206 291454
rect 48970 290898 49206 291134
rect 79690 291218 79926 291454
rect 79690 290898 79926 291134
rect 110410 291218 110646 291454
rect 110410 290898 110646 291134
rect 141130 291218 141366 291454
rect 141130 290898 141366 291134
rect 171850 291218 172086 291454
rect 171850 290898 172086 291134
rect 202570 291218 202806 291454
rect 202570 290898 202806 291134
rect 233290 291218 233526 291454
rect 233290 290898 233526 291134
rect 264010 291218 264246 291454
rect 264010 290898 264246 291134
rect 294730 291218 294966 291454
rect 294730 290898 294966 291134
rect 325450 291218 325686 291454
rect 325450 290898 325686 291134
rect 356170 291218 356406 291454
rect 356170 290898 356406 291134
rect 386890 291218 387126 291454
rect 386890 290898 387126 291134
rect 417610 291218 417846 291454
rect 417610 290898 417846 291134
rect 448330 291218 448566 291454
rect 448330 290898 448566 291134
rect 479050 291218 479286 291454
rect 479050 290898 479286 291134
rect 509770 291218 510006 291454
rect 509770 290898 510006 291134
rect 33610 273218 33846 273454
rect 33610 272898 33846 273134
rect 64330 273218 64566 273454
rect 64330 272898 64566 273134
rect 95050 273218 95286 273454
rect 95050 272898 95286 273134
rect 125770 273218 126006 273454
rect 125770 272898 126006 273134
rect 156490 273218 156726 273454
rect 156490 272898 156726 273134
rect 187210 273218 187446 273454
rect 187210 272898 187446 273134
rect 217930 273218 218166 273454
rect 217930 272898 218166 273134
rect 248650 273218 248886 273454
rect 248650 272898 248886 273134
rect 279370 273218 279606 273454
rect 279370 272898 279606 273134
rect 310090 273218 310326 273454
rect 310090 272898 310326 273134
rect 340810 273218 341046 273454
rect 340810 272898 341046 273134
rect 371530 273218 371766 273454
rect 371530 272898 371766 273134
rect 402250 273218 402486 273454
rect 402250 272898 402486 273134
rect 432970 273218 433206 273454
rect 432970 272898 433206 273134
rect 463690 273218 463926 273454
rect 463690 272898 463926 273134
rect 494410 273218 494646 273454
rect 494410 272898 494646 273134
rect 525130 273218 525366 273454
rect 525130 272898 525366 273134
rect 48970 255218 49206 255454
rect 48970 254898 49206 255134
rect 79690 255218 79926 255454
rect 79690 254898 79926 255134
rect 110410 255218 110646 255454
rect 110410 254898 110646 255134
rect 141130 255218 141366 255454
rect 141130 254898 141366 255134
rect 171850 255218 172086 255454
rect 171850 254898 172086 255134
rect 202570 255218 202806 255454
rect 202570 254898 202806 255134
rect 233290 255218 233526 255454
rect 233290 254898 233526 255134
rect 264010 255218 264246 255454
rect 264010 254898 264246 255134
rect 294730 255218 294966 255454
rect 294730 254898 294966 255134
rect 325450 255218 325686 255454
rect 325450 254898 325686 255134
rect 356170 255218 356406 255454
rect 356170 254898 356406 255134
rect 386890 255218 387126 255454
rect 386890 254898 387126 255134
rect 417610 255218 417846 255454
rect 417610 254898 417846 255134
rect 448330 255218 448566 255454
rect 448330 254898 448566 255134
rect 479050 255218 479286 255454
rect 479050 254898 479286 255134
rect 509770 255218 510006 255454
rect 509770 254898 510006 255134
rect 33610 237218 33846 237454
rect 33610 236898 33846 237134
rect 64330 237218 64566 237454
rect 64330 236898 64566 237134
rect 95050 237218 95286 237454
rect 95050 236898 95286 237134
rect 125770 237218 126006 237454
rect 125770 236898 126006 237134
rect 156490 237218 156726 237454
rect 156490 236898 156726 237134
rect 187210 237218 187446 237454
rect 187210 236898 187446 237134
rect 217930 237218 218166 237454
rect 217930 236898 218166 237134
rect 248650 237218 248886 237454
rect 248650 236898 248886 237134
rect 279370 237218 279606 237454
rect 279370 236898 279606 237134
rect 310090 237218 310326 237454
rect 310090 236898 310326 237134
rect 340810 237218 341046 237454
rect 340810 236898 341046 237134
rect 371530 237218 371766 237454
rect 371530 236898 371766 237134
rect 402250 237218 402486 237454
rect 402250 236898 402486 237134
rect 432970 237218 433206 237454
rect 432970 236898 433206 237134
rect 463690 237218 463926 237454
rect 463690 236898 463926 237134
rect 494410 237218 494646 237454
rect 494410 236898 494646 237134
rect 525130 237218 525366 237454
rect 525130 236898 525366 237134
rect 48970 219218 49206 219454
rect 48970 218898 49206 219134
rect 79690 219218 79926 219454
rect 79690 218898 79926 219134
rect 110410 219218 110646 219454
rect 110410 218898 110646 219134
rect 141130 219218 141366 219454
rect 141130 218898 141366 219134
rect 171850 219218 172086 219454
rect 171850 218898 172086 219134
rect 202570 219218 202806 219454
rect 202570 218898 202806 219134
rect 233290 219218 233526 219454
rect 233290 218898 233526 219134
rect 264010 219218 264246 219454
rect 264010 218898 264246 219134
rect 294730 219218 294966 219454
rect 294730 218898 294966 219134
rect 325450 219218 325686 219454
rect 325450 218898 325686 219134
rect 356170 219218 356406 219454
rect 356170 218898 356406 219134
rect 386890 219218 387126 219454
rect 386890 218898 387126 219134
rect 417610 219218 417846 219454
rect 417610 218898 417846 219134
rect 448330 219218 448566 219454
rect 448330 218898 448566 219134
rect 479050 219218 479286 219454
rect 479050 218898 479286 219134
rect 509770 219218 510006 219454
rect 509770 218898 510006 219134
rect 33610 201218 33846 201454
rect 33610 200898 33846 201134
rect 64330 201218 64566 201454
rect 64330 200898 64566 201134
rect 95050 201218 95286 201454
rect 95050 200898 95286 201134
rect 125770 201218 126006 201454
rect 125770 200898 126006 201134
rect 156490 201218 156726 201454
rect 156490 200898 156726 201134
rect 187210 201218 187446 201454
rect 187210 200898 187446 201134
rect 217930 201218 218166 201454
rect 217930 200898 218166 201134
rect 248650 201218 248886 201454
rect 248650 200898 248886 201134
rect 279370 201218 279606 201454
rect 279370 200898 279606 201134
rect 310090 201218 310326 201454
rect 310090 200898 310326 201134
rect 340810 201218 341046 201454
rect 340810 200898 341046 201134
rect 371530 201218 371766 201454
rect 371530 200898 371766 201134
rect 402250 201218 402486 201454
rect 402250 200898 402486 201134
rect 432970 201218 433206 201454
rect 432970 200898 433206 201134
rect 463690 201218 463926 201454
rect 463690 200898 463926 201134
rect 494410 201218 494646 201454
rect 494410 200898 494646 201134
rect 525130 201218 525366 201454
rect 525130 200898 525366 201134
rect 48970 183218 49206 183454
rect 48970 182898 49206 183134
rect 79690 183218 79926 183454
rect 79690 182898 79926 183134
rect 110410 183218 110646 183454
rect 110410 182898 110646 183134
rect 141130 183218 141366 183454
rect 141130 182898 141366 183134
rect 171850 183218 172086 183454
rect 171850 182898 172086 183134
rect 202570 183218 202806 183454
rect 202570 182898 202806 183134
rect 233290 183218 233526 183454
rect 233290 182898 233526 183134
rect 264010 183218 264246 183454
rect 264010 182898 264246 183134
rect 294730 183218 294966 183454
rect 294730 182898 294966 183134
rect 325450 183218 325686 183454
rect 325450 182898 325686 183134
rect 356170 183218 356406 183454
rect 356170 182898 356406 183134
rect 386890 183218 387126 183454
rect 386890 182898 387126 183134
rect 417610 183218 417846 183454
rect 417610 182898 417846 183134
rect 448330 183218 448566 183454
rect 448330 182898 448566 183134
rect 479050 183218 479286 183454
rect 479050 182898 479286 183134
rect 509770 183218 510006 183454
rect 509770 182898 510006 183134
rect 33610 165218 33846 165454
rect 33610 164898 33846 165134
rect 64330 165218 64566 165454
rect 64330 164898 64566 165134
rect 95050 165218 95286 165454
rect 95050 164898 95286 165134
rect 125770 165218 126006 165454
rect 125770 164898 126006 165134
rect 156490 165218 156726 165454
rect 156490 164898 156726 165134
rect 187210 165218 187446 165454
rect 187210 164898 187446 165134
rect 217930 165218 218166 165454
rect 217930 164898 218166 165134
rect 248650 165218 248886 165454
rect 248650 164898 248886 165134
rect 279370 165218 279606 165454
rect 279370 164898 279606 165134
rect 310090 165218 310326 165454
rect 310090 164898 310326 165134
rect 340810 165218 341046 165454
rect 340810 164898 341046 165134
rect 371530 165218 371766 165454
rect 371530 164898 371766 165134
rect 402250 165218 402486 165454
rect 402250 164898 402486 165134
rect 432970 165218 433206 165454
rect 432970 164898 433206 165134
rect 463690 165218 463926 165454
rect 463690 164898 463926 165134
rect 494410 165218 494646 165454
rect 494410 164898 494646 165134
rect 525130 165218 525366 165454
rect 525130 164898 525366 165134
rect 48970 147218 49206 147454
rect 48970 146898 49206 147134
rect 79690 147218 79926 147454
rect 79690 146898 79926 147134
rect 110410 147218 110646 147454
rect 110410 146898 110646 147134
rect 141130 147218 141366 147454
rect 141130 146898 141366 147134
rect 171850 147218 172086 147454
rect 171850 146898 172086 147134
rect 202570 147218 202806 147454
rect 202570 146898 202806 147134
rect 233290 147218 233526 147454
rect 233290 146898 233526 147134
rect 264010 147218 264246 147454
rect 264010 146898 264246 147134
rect 294730 147218 294966 147454
rect 294730 146898 294966 147134
rect 325450 147218 325686 147454
rect 325450 146898 325686 147134
rect 356170 147218 356406 147454
rect 356170 146898 356406 147134
rect 386890 147218 387126 147454
rect 386890 146898 387126 147134
rect 417610 147218 417846 147454
rect 417610 146898 417846 147134
rect 448330 147218 448566 147454
rect 448330 146898 448566 147134
rect 479050 147218 479286 147454
rect 479050 146898 479286 147134
rect 509770 147218 510006 147454
rect 509770 146898 510006 147134
rect 33610 129218 33846 129454
rect 33610 128898 33846 129134
rect 64330 129218 64566 129454
rect 64330 128898 64566 129134
rect 95050 129218 95286 129454
rect 95050 128898 95286 129134
rect 125770 129218 126006 129454
rect 125770 128898 126006 129134
rect 156490 129218 156726 129454
rect 156490 128898 156726 129134
rect 187210 129218 187446 129454
rect 187210 128898 187446 129134
rect 217930 129218 218166 129454
rect 217930 128898 218166 129134
rect 248650 129218 248886 129454
rect 248650 128898 248886 129134
rect 279370 129218 279606 129454
rect 279370 128898 279606 129134
rect 310090 129218 310326 129454
rect 310090 128898 310326 129134
rect 340810 129218 341046 129454
rect 340810 128898 341046 129134
rect 371530 129218 371766 129454
rect 371530 128898 371766 129134
rect 402250 129218 402486 129454
rect 402250 128898 402486 129134
rect 432970 129218 433206 129454
rect 432970 128898 433206 129134
rect 463690 129218 463926 129454
rect 463690 128898 463926 129134
rect 494410 129218 494646 129454
rect 494410 128898 494646 129134
rect 525130 129218 525366 129454
rect 525130 128898 525366 129134
rect 48970 111218 49206 111454
rect 48970 110898 49206 111134
rect 79690 111218 79926 111454
rect 79690 110898 79926 111134
rect 110410 111218 110646 111454
rect 110410 110898 110646 111134
rect 141130 111218 141366 111454
rect 141130 110898 141366 111134
rect 171850 111218 172086 111454
rect 171850 110898 172086 111134
rect 202570 111218 202806 111454
rect 202570 110898 202806 111134
rect 233290 111218 233526 111454
rect 233290 110898 233526 111134
rect 264010 111218 264246 111454
rect 264010 110898 264246 111134
rect 294730 111218 294966 111454
rect 294730 110898 294966 111134
rect 325450 111218 325686 111454
rect 325450 110898 325686 111134
rect 356170 111218 356406 111454
rect 356170 110898 356406 111134
rect 386890 111218 387126 111454
rect 386890 110898 387126 111134
rect 417610 111218 417846 111454
rect 417610 110898 417846 111134
rect 448330 111218 448566 111454
rect 448330 110898 448566 111134
rect 479050 111218 479286 111454
rect 479050 110898 479286 111134
rect 509770 111218 510006 111454
rect 509770 110898 510006 111134
rect 33610 93218 33846 93454
rect 33610 92898 33846 93134
rect 64330 93218 64566 93454
rect 64330 92898 64566 93134
rect 95050 93218 95286 93454
rect 95050 92898 95286 93134
rect 125770 93218 126006 93454
rect 125770 92898 126006 93134
rect 156490 93218 156726 93454
rect 156490 92898 156726 93134
rect 187210 93218 187446 93454
rect 187210 92898 187446 93134
rect 217930 93218 218166 93454
rect 217930 92898 218166 93134
rect 248650 93218 248886 93454
rect 248650 92898 248886 93134
rect 279370 93218 279606 93454
rect 279370 92898 279606 93134
rect 310090 93218 310326 93454
rect 310090 92898 310326 93134
rect 340810 93218 341046 93454
rect 340810 92898 341046 93134
rect 371530 93218 371766 93454
rect 371530 92898 371766 93134
rect 402250 93218 402486 93454
rect 402250 92898 402486 93134
rect 432970 93218 433206 93454
rect 432970 92898 433206 93134
rect 463690 93218 463926 93454
rect 463690 92898 463926 93134
rect 494410 93218 494646 93454
rect 494410 92898 494646 93134
rect 525130 93218 525366 93454
rect 525130 92898 525366 93134
rect 48970 75218 49206 75454
rect 48970 74898 49206 75134
rect 79690 75218 79926 75454
rect 79690 74898 79926 75134
rect 110410 75218 110646 75454
rect 110410 74898 110646 75134
rect 141130 75218 141366 75454
rect 141130 74898 141366 75134
rect 171850 75218 172086 75454
rect 171850 74898 172086 75134
rect 202570 75218 202806 75454
rect 202570 74898 202806 75134
rect 233290 75218 233526 75454
rect 233290 74898 233526 75134
rect 264010 75218 264246 75454
rect 264010 74898 264246 75134
rect 294730 75218 294966 75454
rect 294730 74898 294966 75134
rect 325450 75218 325686 75454
rect 325450 74898 325686 75134
rect 356170 75218 356406 75454
rect 356170 74898 356406 75134
rect 386890 75218 387126 75454
rect 386890 74898 387126 75134
rect 417610 75218 417846 75454
rect 417610 74898 417846 75134
rect 448330 75218 448566 75454
rect 448330 74898 448566 75134
rect 479050 75218 479286 75454
rect 479050 74898 479286 75134
rect 509770 75218 510006 75454
rect 509770 74898 510006 75134
rect 33610 57218 33846 57454
rect 33610 56898 33846 57134
rect 64330 57218 64566 57454
rect 64330 56898 64566 57134
rect 95050 57218 95286 57454
rect 95050 56898 95286 57134
rect 125770 57218 126006 57454
rect 125770 56898 126006 57134
rect 156490 57218 156726 57454
rect 156490 56898 156726 57134
rect 187210 57218 187446 57454
rect 187210 56898 187446 57134
rect 217930 57218 218166 57454
rect 217930 56898 218166 57134
rect 248650 57218 248886 57454
rect 248650 56898 248886 57134
rect 279370 57218 279606 57454
rect 279370 56898 279606 57134
rect 310090 57218 310326 57454
rect 310090 56898 310326 57134
rect 340810 57218 341046 57454
rect 340810 56898 341046 57134
rect 371530 57218 371766 57454
rect 371530 56898 371766 57134
rect 402250 57218 402486 57454
rect 402250 56898 402486 57134
rect 432970 57218 433206 57454
rect 432970 56898 433206 57134
rect 463690 57218 463926 57454
rect 463690 56898 463926 57134
rect 494410 57218 494646 57454
rect 494410 56898 494646 57134
rect 525130 57218 525366 57454
rect 525130 56898 525366 57134
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 540490 651218 540726 651454
rect 540490 650898 540726 651134
rect 540490 615218 540726 615454
rect 540490 614898 540726 615134
rect 540490 579218 540726 579454
rect 540490 578898 540726 579134
rect 540490 543218 540726 543454
rect 540490 542898 540726 543134
rect 540490 507218 540726 507454
rect 540490 506898 540726 507134
rect 540014 484382 540250 484618
rect 540934 484532 541170 484618
rect 540934 484468 541020 484532
rect 541020 484468 541084 484532
rect 541084 484468 541170 484532
rect 540934 484382 541170 484468
rect 540490 471218 540726 471454
rect 540490 470898 540726 471134
rect 540490 435218 540726 435454
rect 540490 434898 540726 435134
rect 540490 399218 540726 399454
rect 540490 398898 540726 399134
rect 540490 363218 540726 363454
rect 540490 362898 540726 363134
rect 540490 327218 540726 327454
rect 540490 326898 540726 327134
rect 540490 291218 540726 291454
rect 540490 290898 540726 291134
rect 540490 255218 540726 255454
rect 540490 254898 540726 255134
rect 540490 219218 540726 219454
rect 540490 218898 540726 219134
rect 540490 183218 540726 183454
rect 540490 182898 540726 183134
rect 540490 147218 540726 147454
rect 540490 146898 540726 147134
rect 540490 111218 540726 111454
rect 540490 110898 540726 111134
rect 540490 75218 540726 75454
rect 540490 74898 540726 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 18250 651454
rect 18486 651218 48970 651454
rect 49206 651218 79690 651454
rect 79926 651218 110410 651454
rect 110646 651218 141130 651454
rect 141366 651218 171850 651454
rect 172086 651218 202570 651454
rect 202806 651218 233290 651454
rect 233526 651218 264010 651454
rect 264246 651218 294730 651454
rect 294966 651218 325450 651454
rect 325686 651218 356170 651454
rect 356406 651218 386890 651454
rect 387126 651218 417610 651454
rect 417846 651218 448330 651454
rect 448566 651218 479050 651454
rect 479286 651218 509770 651454
rect 510006 651218 540490 651454
rect 540726 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 18250 651134
rect 18486 650898 48970 651134
rect 49206 650898 79690 651134
rect 79926 650898 110410 651134
rect 110646 650898 141130 651134
rect 141366 650898 171850 651134
rect 172086 650898 202570 651134
rect 202806 650898 233290 651134
rect 233526 650898 264010 651134
rect 264246 650898 294730 651134
rect 294966 650898 325450 651134
rect 325686 650898 356170 651134
rect 356406 650898 386890 651134
rect 387126 650898 417610 651134
rect 417846 650898 448330 651134
rect 448566 650898 479050 651134
rect 479286 650898 509770 651134
rect 510006 650898 540490 651134
rect 540726 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 33610 633454
rect 33846 633218 64330 633454
rect 64566 633218 95050 633454
rect 95286 633218 125770 633454
rect 126006 633218 156490 633454
rect 156726 633218 187210 633454
rect 187446 633218 217930 633454
rect 218166 633218 248650 633454
rect 248886 633218 279370 633454
rect 279606 633218 310090 633454
rect 310326 633218 340810 633454
rect 341046 633218 371530 633454
rect 371766 633218 402250 633454
rect 402486 633218 432970 633454
rect 433206 633218 463690 633454
rect 463926 633218 494410 633454
rect 494646 633218 525130 633454
rect 525366 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 33610 633134
rect 33846 632898 64330 633134
rect 64566 632898 95050 633134
rect 95286 632898 125770 633134
rect 126006 632898 156490 633134
rect 156726 632898 187210 633134
rect 187446 632898 217930 633134
rect 218166 632898 248650 633134
rect 248886 632898 279370 633134
rect 279606 632898 310090 633134
rect 310326 632898 340810 633134
rect 341046 632898 371530 633134
rect 371766 632898 402250 633134
rect 402486 632898 432970 633134
rect 433206 632898 463690 633134
rect 463926 632898 494410 633134
rect 494646 632898 525130 633134
rect 525366 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 18250 615454
rect 18486 615218 48970 615454
rect 49206 615218 79690 615454
rect 79926 615218 110410 615454
rect 110646 615218 141130 615454
rect 141366 615218 171850 615454
rect 172086 615218 202570 615454
rect 202806 615218 233290 615454
rect 233526 615218 264010 615454
rect 264246 615218 294730 615454
rect 294966 615218 325450 615454
rect 325686 615218 356170 615454
rect 356406 615218 386890 615454
rect 387126 615218 417610 615454
rect 417846 615218 448330 615454
rect 448566 615218 479050 615454
rect 479286 615218 509770 615454
rect 510006 615218 540490 615454
rect 540726 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 18250 615134
rect 18486 614898 48970 615134
rect 49206 614898 79690 615134
rect 79926 614898 110410 615134
rect 110646 614898 141130 615134
rect 141366 614898 171850 615134
rect 172086 614898 202570 615134
rect 202806 614898 233290 615134
rect 233526 614898 264010 615134
rect 264246 614898 294730 615134
rect 294966 614898 325450 615134
rect 325686 614898 356170 615134
rect 356406 614898 386890 615134
rect 387126 614898 417610 615134
rect 417846 614898 448330 615134
rect 448566 614898 479050 615134
rect 479286 614898 509770 615134
rect 510006 614898 540490 615134
rect 540726 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 33610 597454
rect 33846 597218 64330 597454
rect 64566 597218 95050 597454
rect 95286 597218 125770 597454
rect 126006 597218 156490 597454
rect 156726 597218 187210 597454
rect 187446 597218 217930 597454
rect 218166 597218 248650 597454
rect 248886 597218 279370 597454
rect 279606 597218 310090 597454
rect 310326 597218 340810 597454
rect 341046 597218 371530 597454
rect 371766 597218 402250 597454
rect 402486 597218 432970 597454
rect 433206 597218 463690 597454
rect 463926 597218 494410 597454
rect 494646 597218 525130 597454
rect 525366 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 33610 597134
rect 33846 596898 64330 597134
rect 64566 596898 95050 597134
rect 95286 596898 125770 597134
rect 126006 596898 156490 597134
rect 156726 596898 187210 597134
rect 187446 596898 217930 597134
rect 218166 596898 248650 597134
rect 248886 596898 279370 597134
rect 279606 596898 310090 597134
rect 310326 596898 340810 597134
rect 341046 596898 371530 597134
rect 371766 596898 402250 597134
rect 402486 596898 432970 597134
rect 433206 596898 463690 597134
rect 463926 596898 494410 597134
rect 494646 596898 525130 597134
rect 525366 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 18250 579454
rect 18486 579218 48970 579454
rect 49206 579218 79690 579454
rect 79926 579218 110410 579454
rect 110646 579218 141130 579454
rect 141366 579218 171850 579454
rect 172086 579218 202570 579454
rect 202806 579218 233290 579454
rect 233526 579218 264010 579454
rect 264246 579218 294730 579454
rect 294966 579218 325450 579454
rect 325686 579218 356170 579454
rect 356406 579218 386890 579454
rect 387126 579218 417610 579454
rect 417846 579218 448330 579454
rect 448566 579218 479050 579454
rect 479286 579218 509770 579454
rect 510006 579218 540490 579454
rect 540726 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 18250 579134
rect 18486 578898 48970 579134
rect 49206 578898 79690 579134
rect 79926 578898 110410 579134
rect 110646 578898 141130 579134
rect 141366 578898 171850 579134
rect 172086 578898 202570 579134
rect 202806 578898 233290 579134
rect 233526 578898 264010 579134
rect 264246 578898 294730 579134
rect 294966 578898 325450 579134
rect 325686 578898 356170 579134
rect 356406 578898 386890 579134
rect 387126 578898 417610 579134
rect 417846 578898 448330 579134
rect 448566 578898 479050 579134
rect 479286 578898 509770 579134
rect 510006 578898 540490 579134
rect 540726 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 33610 561454
rect 33846 561218 64330 561454
rect 64566 561218 95050 561454
rect 95286 561218 125770 561454
rect 126006 561218 156490 561454
rect 156726 561218 187210 561454
rect 187446 561218 217930 561454
rect 218166 561218 248650 561454
rect 248886 561218 279370 561454
rect 279606 561218 310090 561454
rect 310326 561218 340810 561454
rect 341046 561218 371530 561454
rect 371766 561218 402250 561454
rect 402486 561218 432970 561454
rect 433206 561218 463690 561454
rect 463926 561218 494410 561454
rect 494646 561218 525130 561454
rect 525366 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 33610 561134
rect 33846 560898 64330 561134
rect 64566 560898 95050 561134
rect 95286 560898 125770 561134
rect 126006 560898 156490 561134
rect 156726 560898 187210 561134
rect 187446 560898 217930 561134
rect 218166 560898 248650 561134
rect 248886 560898 279370 561134
rect 279606 560898 310090 561134
rect 310326 560898 340810 561134
rect 341046 560898 371530 561134
rect 371766 560898 402250 561134
rect 402486 560898 432970 561134
rect 433206 560898 463690 561134
rect 463926 560898 494410 561134
rect 494646 560898 525130 561134
rect 525366 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 18250 543454
rect 18486 543218 48970 543454
rect 49206 543218 79690 543454
rect 79926 543218 110410 543454
rect 110646 543218 141130 543454
rect 141366 543218 171850 543454
rect 172086 543218 202570 543454
rect 202806 543218 233290 543454
rect 233526 543218 264010 543454
rect 264246 543218 294730 543454
rect 294966 543218 325450 543454
rect 325686 543218 356170 543454
rect 356406 543218 386890 543454
rect 387126 543218 417610 543454
rect 417846 543218 448330 543454
rect 448566 543218 479050 543454
rect 479286 543218 509770 543454
rect 510006 543218 540490 543454
rect 540726 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 18250 543134
rect 18486 542898 48970 543134
rect 49206 542898 79690 543134
rect 79926 542898 110410 543134
rect 110646 542898 141130 543134
rect 141366 542898 171850 543134
rect 172086 542898 202570 543134
rect 202806 542898 233290 543134
rect 233526 542898 264010 543134
rect 264246 542898 294730 543134
rect 294966 542898 325450 543134
rect 325686 542898 356170 543134
rect 356406 542898 386890 543134
rect 387126 542898 417610 543134
rect 417846 542898 448330 543134
rect 448566 542898 479050 543134
rect 479286 542898 509770 543134
rect 510006 542898 540490 543134
rect 540726 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 33610 525454
rect 33846 525218 64330 525454
rect 64566 525218 95050 525454
rect 95286 525218 125770 525454
rect 126006 525218 156490 525454
rect 156726 525218 187210 525454
rect 187446 525218 217930 525454
rect 218166 525218 248650 525454
rect 248886 525218 279370 525454
rect 279606 525218 310090 525454
rect 310326 525218 340810 525454
rect 341046 525218 371530 525454
rect 371766 525218 402250 525454
rect 402486 525218 432970 525454
rect 433206 525218 463690 525454
rect 463926 525218 494410 525454
rect 494646 525218 525130 525454
rect 525366 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 33610 525134
rect 33846 524898 64330 525134
rect 64566 524898 95050 525134
rect 95286 524898 125770 525134
rect 126006 524898 156490 525134
rect 156726 524898 187210 525134
rect 187446 524898 217930 525134
rect 218166 524898 248650 525134
rect 248886 524898 279370 525134
rect 279606 524898 310090 525134
rect 310326 524898 340810 525134
rect 341046 524898 371530 525134
rect 371766 524898 402250 525134
rect 402486 524898 432970 525134
rect 433206 524898 463690 525134
rect 463926 524898 494410 525134
rect 494646 524898 525130 525134
rect 525366 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 18250 507454
rect 18486 507218 48970 507454
rect 49206 507218 79690 507454
rect 79926 507218 110410 507454
rect 110646 507218 141130 507454
rect 141366 507218 171850 507454
rect 172086 507218 202570 507454
rect 202806 507218 233290 507454
rect 233526 507218 264010 507454
rect 264246 507218 294730 507454
rect 294966 507218 325450 507454
rect 325686 507218 356170 507454
rect 356406 507218 386890 507454
rect 387126 507218 417610 507454
rect 417846 507218 448330 507454
rect 448566 507218 479050 507454
rect 479286 507218 509770 507454
rect 510006 507218 540490 507454
rect 540726 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 18250 507134
rect 18486 506898 48970 507134
rect 49206 506898 79690 507134
rect 79926 506898 110410 507134
rect 110646 506898 141130 507134
rect 141366 506898 171850 507134
rect 172086 506898 202570 507134
rect 202806 506898 233290 507134
rect 233526 506898 264010 507134
rect 264246 506898 294730 507134
rect 294966 506898 325450 507134
rect 325686 506898 356170 507134
rect 356406 506898 386890 507134
rect 387126 506898 417610 507134
rect 417846 506898 448330 507134
rect 448566 506898 479050 507134
rect 479286 506898 509770 507134
rect 510006 506898 540490 507134
rect 540726 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 33610 489454
rect 33846 489218 64330 489454
rect 64566 489218 95050 489454
rect 95286 489218 125770 489454
rect 126006 489218 156490 489454
rect 156726 489218 187210 489454
rect 187446 489218 217930 489454
rect 218166 489218 248650 489454
rect 248886 489218 279370 489454
rect 279606 489218 310090 489454
rect 310326 489218 340810 489454
rect 341046 489218 371530 489454
rect 371766 489218 402250 489454
rect 402486 489218 432970 489454
rect 433206 489218 463690 489454
rect 463926 489218 494410 489454
rect 494646 489218 525130 489454
rect 525366 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 33610 489134
rect 33846 488898 64330 489134
rect 64566 488898 95050 489134
rect 95286 488898 125770 489134
rect 126006 488898 156490 489134
rect 156726 488898 187210 489134
rect 187446 488898 217930 489134
rect 218166 488898 248650 489134
rect 248886 488898 279370 489134
rect 279606 488898 310090 489134
rect 310326 488898 340810 489134
rect 341046 488898 371530 489134
rect 371766 488898 402250 489134
rect 402486 488898 432970 489134
rect 433206 488898 463690 489134
rect 463926 488898 494410 489134
rect 494646 488898 525130 489134
rect 525366 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect 539972 484618 541212 484660
rect 539972 484382 540014 484618
rect 540250 484382 540934 484618
rect 541170 484382 541212 484618
rect 539972 484340 541212 484382
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 18250 471454
rect 18486 471218 48970 471454
rect 49206 471218 79690 471454
rect 79926 471218 110410 471454
rect 110646 471218 141130 471454
rect 141366 471218 171850 471454
rect 172086 471218 202570 471454
rect 202806 471218 233290 471454
rect 233526 471218 264010 471454
rect 264246 471218 294730 471454
rect 294966 471218 325450 471454
rect 325686 471218 356170 471454
rect 356406 471218 386890 471454
rect 387126 471218 417610 471454
rect 417846 471218 448330 471454
rect 448566 471218 479050 471454
rect 479286 471218 509770 471454
rect 510006 471218 540490 471454
rect 540726 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 18250 471134
rect 18486 470898 48970 471134
rect 49206 470898 79690 471134
rect 79926 470898 110410 471134
rect 110646 470898 141130 471134
rect 141366 470898 171850 471134
rect 172086 470898 202570 471134
rect 202806 470898 233290 471134
rect 233526 470898 264010 471134
rect 264246 470898 294730 471134
rect 294966 470898 325450 471134
rect 325686 470898 356170 471134
rect 356406 470898 386890 471134
rect 387126 470898 417610 471134
rect 417846 470898 448330 471134
rect 448566 470898 479050 471134
rect 479286 470898 509770 471134
rect 510006 470898 540490 471134
rect 540726 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 33610 453454
rect 33846 453218 64330 453454
rect 64566 453218 95050 453454
rect 95286 453218 125770 453454
rect 126006 453218 156490 453454
rect 156726 453218 187210 453454
rect 187446 453218 217930 453454
rect 218166 453218 248650 453454
rect 248886 453218 279370 453454
rect 279606 453218 310090 453454
rect 310326 453218 340810 453454
rect 341046 453218 371530 453454
rect 371766 453218 402250 453454
rect 402486 453218 432970 453454
rect 433206 453218 463690 453454
rect 463926 453218 494410 453454
rect 494646 453218 525130 453454
rect 525366 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 33610 453134
rect 33846 452898 64330 453134
rect 64566 452898 95050 453134
rect 95286 452898 125770 453134
rect 126006 452898 156490 453134
rect 156726 452898 187210 453134
rect 187446 452898 217930 453134
rect 218166 452898 248650 453134
rect 248886 452898 279370 453134
rect 279606 452898 310090 453134
rect 310326 452898 340810 453134
rect 341046 452898 371530 453134
rect 371766 452898 402250 453134
rect 402486 452898 432970 453134
rect 433206 452898 463690 453134
rect 463926 452898 494410 453134
rect 494646 452898 525130 453134
rect 525366 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 18250 435454
rect 18486 435218 48970 435454
rect 49206 435218 79690 435454
rect 79926 435218 110410 435454
rect 110646 435218 141130 435454
rect 141366 435218 171850 435454
rect 172086 435218 202570 435454
rect 202806 435218 233290 435454
rect 233526 435218 264010 435454
rect 264246 435218 294730 435454
rect 294966 435218 325450 435454
rect 325686 435218 356170 435454
rect 356406 435218 386890 435454
rect 387126 435218 417610 435454
rect 417846 435218 448330 435454
rect 448566 435218 479050 435454
rect 479286 435218 509770 435454
rect 510006 435218 540490 435454
rect 540726 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 18250 435134
rect 18486 434898 48970 435134
rect 49206 434898 79690 435134
rect 79926 434898 110410 435134
rect 110646 434898 141130 435134
rect 141366 434898 171850 435134
rect 172086 434898 202570 435134
rect 202806 434898 233290 435134
rect 233526 434898 264010 435134
rect 264246 434898 294730 435134
rect 294966 434898 325450 435134
rect 325686 434898 356170 435134
rect 356406 434898 386890 435134
rect 387126 434898 417610 435134
rect 417846 434898 448330 435134
rect 448566 434898 479050 435134
rect 479286 434898 509770 435134
rect 510006 434898 540490 435134
rect 540726 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 33610 417454
rect 33846 417218 64330 417454
rect 64566 417218 95050 417454
rect 95286 417218 125770 417454
rect 126006 417218 156490 417454
rect 156726 417218 187210 417454
rect 187446 417218 217930 417454
rect 218166 417218 248650 417454
rect 248886 417218 279370 417454
rect 279606 417218 310090 417454
rect 310326 417218 340810 417454
rect 341046 417218 371530 417454
rect 371766 417218 402250 417454
rect 402486 417218 432970 417454
rect 433206 417218 463690 417454
rect 463926 417218 494410 417454
rect 494646 417218 525130 417454
rect 525366 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 33610 417134
rect 33846 416898 64330 417134
rect 64566 416898 95050 417134
rect 95286 416898 125770 417134
rect 126006 416898 156490 417134
rect 156726 416898 187210 417134
rect 187446 416898 217930 417134
rect 218166 416898 248650 417134
rect 248886 416898 279370 417134
rect 279606 416898 310090 417134
rect 310326 416898 340810 417134
rect 341046 416898 371530 417134
rect 371766 416898 402250 417134
rect 402486 416898 432970 417134
rect 433206 416898 463690 417134
rect 463926 416898 494410 417134
rect 494646 416898 525130 417134
rect 525366 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 18250 399454
rect 18486 399218 48970 399454
rect 49206 399218 79690 399454
rect 79926 399218 110410 399454
rect 110646 399218 141130 399454
rect 141366 399218 171850 399454
rect 172086 399218 202570 399454
rect 202806 399218 233290 399454
rect 233526 399218 264010 399454
rect 264246 399218 294730 399454
rect 294966 399218 325450 399454
rect 325686 399218 356170 399454
rect 356406 399218 386890 399454
rect 387126 399218 417610 399454
rect 417846 399218 448330 399454
rect 448566 399218 479050 399454
rect 479286 399218 509770 399454
rect 510006 399218 540490 399454
rect 540726 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 18250 399134
rect 18486 398898 48970 399134
rect 49206 398898 79690 399134
rect 79926 398898 110410 399134
rect 110646 398898 141130 399134
rect 141366 398898 171850 399134
rect 172086 398898 202570 399134
rect 202806 398898 233290 399134
rect 233526 398898 264010 399134
rect 264246 398898 294730 399134
rect 294966 398898 325450 399134
rect 325686 398898 356170 399134
rect 356406 398898 386890 399134
rect 387126 398898 417610 399134
rect 417846 398898 448330 399134
rect 448566 398898 479050 399134
rect 479286 398898 509770 399134
rect 510006 398898 540490 399134
rect 540726 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 33610 381454
rect 33846 381218 64330 381454
rect 64566 381218 95050 381454
rect 95286 381218 125770 381454
rect 126006 381218 156490 381454
rect 156726 381218 187210 381454
rect 187446 381218 217930 381454
rect 218166 381218 248650 381454
rect 248886 381218 279370 381454
rect 279606 381218 310090 381454
rect 310326 381218 340810 381454
rect 341046 381218 371530 381454
rect 371766 381218 402250 381454
rect 402486 381218 432970 381454
rect 433206 381218 463690 381454
rect 463926 381218 494410 381454
rect 494646 381218 525130 381454
rect 525366 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 33610 381134
rect 33846 380898 64330 381134
rect 64566 380898 95050 381134
rect 95286 380898 125770 381134
rect 126006 380898 156490 381134
rect 156726 380898 187210 381134
rect 187446 380898 217930 381134
rect 218166 380898 248650 381134
rect 248886 380898 279370 381134
rect 279606 380898 310090 381134
rect 310326 380898 340810 381134
rect 341046 380898 371530 381134
rect 371766 380898 402250 381134
rect 402486 380898 432970 381134
rect 433206 380898 463690 381134
rect 463926 380898 494410 381134
rect 494646 380898 525130 381134
rect 525366 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 18250 363454
rect 18486 363218 48970 363454
rect 49206 363218 79690 363454
rect 79926 363218 110410 363454
rect 110646 363218 141130 363454
rect 141366 363218 171850 363454
rect 172086 363218 202570 363454
rect 202806 363218 233290 363454
rect 233526 363218 264010 363454
rect 264246 363218 294730 363454
rect 294966 363218 325450 363454
rect 325686 363218 356170 363454
rect 356406 363218 386890 363454
rect 387126 363218 417610 363454
rect 417846 363218 448330 363454
rect 448566 363218 479050 363454
rect 479286 363218 509770 363454
rect 510006 363218 540490 363454
rect 540726 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 18250 363134
rect 18486 362898 48970 363134
rect 49206 362898 79690 363134
rect 79926 362898 110410 363134
rect 110646 362898 141130 363134
rect 141366 362898 171850 363134
rect 172086 362898 202570 363134
rect 202806 362898 233290 363134
rect 233526 362898 264010 363134
rect 264246 362898 294730 363134
rect 294966 362898 325450 363134
rect 325686 362898 356170 363134
rect 356406 362898 386890 363134
rect 387126 362898 417610 363134
rect 417846 362898 448330 363134
rect 448566 362898 479050 363134
rect 479286 362898 509770 363134
rect 510006 362898 540490 363134
rect 540726 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 33610 345454
rect 33846 345218 64330 345454
rect 64566 345218 95050 345454
rect 95286 345218 125770 345454
rect 126006 345218 156490 345454
rect 156726 345218 187210 345454
rect 187446 345218 217930 345454
rect 218166 345218 248650 345454
rect 248886 345218 279370 345454
rect 279606 345218 310090 345454
rect 310326 345218 340810 345454
rect 341046 345218 371530 345454
rect 371766 345218 402250 345454
rect 402486 345218 432970 345454
rect 433206 345218 463690 345454
rect 463926 345218 494410 345454
rect 494646 345218 525130 345454
rect 525366 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 33610 345134
rect 33846 344898 64330 345134
rect 64566 344898 95050 345134
rect 95286 344898 125770 345134
rect 126006 344898 156490 345134
rect 156726 344898 187210 345134
rect 187446 344898 217930 345134
rect 218166 344898 248650 345134
rect 248886 344898 279370 345134
rect 279606 344898 310090 345134
rect 310326 344898 340810 345134
rect 341046 344898 371530 345134
rect 371766 344898 402250 345134
rect 402486 344898 432970 345134
rect 433206 344898 463690 345134
rect 463926 344898 494410 345134
rect 494646 344898 525130 345134
rect 525366 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 18250 327454
rect 18486 327218 48970 327454
rect 49206 327218 79690 327454
rect 79926 327218 110410 327454
rect 110646 327218 141130 327454
rect 141366 327218 171850 327454
rect 172086 327218 202570 327454
rect 202806 327218 233290 327454
rect 233526 327218 264010 327454
rect 264246 327218 294730 327454
rect 294966 327218 325450 327454
rect 325686 327218 356170 327454
rect 356406 327218 386890 327454
rect 387126 327218 417610 327454
rect 417846 327218 448330 327454
rect 448566 327218 479050 327454
rect 479286 327218 509770 327454
rect 510006 327218 540490 327454
rect 540726 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 18250 327134
rect 18486 326898 48970 327134
rect 49206 326898 79690 327134
rect 79926 326898 110410 327134
rect 110646 326898 141130 327134
rect 141366 326898 171850 327134
rect 172086 326898 202570 327134
rect 202806 326898 233290 327134
rect 233526 326898 264010 327134
rect 264246 326898 294730 327134
rect 294966 326898 325450 327134
rect 325686 326898 356170 327134
rect 356406 326898 386890 327134
rect 387126 326898 417610 327134
rect 417846 326898 448330 327134
rect 448566 326898 479050 327134
rect 479286 326898 509770 327134
rect 510006 326898 540490 327134
rect 540726 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 33610 309454
rect 33846 309218 64330 309454
rect 64566 309218 95050 309454
rect 95286 309218 125770 309454
rect 126006 309218 156490 309454
rect 156726 309218 187210 309454
rect 187446 309218 217930 309454
rect 218166 309218 248650 309454
rect 248886 309218 279370 309454
rect 279606 309218 310090 309454
rect 310326 309218 340810 309454
rect 341046 309218 371530 309454
rect 371766 309218 402250 309454
rect 402486 309218 432970 309454
rect 433206 309218 463690 309454
rect 463926 309218 494410 309454
rect 494646 309218 525130 309454
rect 525366 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 33610 309134
rect 33846 308898 64330 309134
rect 64566 308898 95050 309134
rect 95286 308898 125770 309134
rect 126006 308898 156490 309134
rect 156726 308898 187210 309134
rect 187446 308898 217930 309134
rect 218166 308898 248650 309134
rect 248886 308898 279370 309134
rect 279606 308898 310090 309134
rect 310326 308898 340810 309134
rect 341046 308898 371530 309134
rect 371766 308898 402250 309134
rect 402486 308898 432970 309134
rect 433206 308898 463690 309134
rect 463926 308898 494410 309134
rect 494646 308898 525130 309134
rect 525366 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 18250 291454
rect 18486 291218 48970 291454
rect 49206 291218 79690 291454
rect 79926 291218 110410 291454
rect 110646 291218 141130 291454
rect 141366 291218 171850 291454
rect 172086 291218 202570 291454
rect 202806 291218 233290 291454
rect 233526 291218 264010 291454
rect 264246 291218 294730 291454
rect 294966 291218 325450 291454
rect 325686 291218 356170 291454
rect 356406 291218 386890 291454
rect 387126 291218 417610 291454
rect 417846 291218 448330 291454
rect 448566 291218 479050 291454
rect 479286 291218 509770 291454
rect 510006 291218 540490 291454
rect 540726 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 18250 291134
rect 18486 290898 48970 291134
rect 49206 290898 79690 291134
rect 79926 290898 110410 291134
rect 110646 290898 141130 291134
rect 141366 290898 171850 291134
rect 172086 290898 202570 291134
rect 202806 290898 233290 291134
rect 233526 290898 264010 291134
rect 264246 290898 294730 291134
rect 294966 290898 325450 291134
rect 325686 290898 356170 291134
rect 356406 290898 386890 291134
rect 387126 290898 417610 291134
rect 417846 290898 448330 291134
rect 448566 290898 479050 291134
rect 479286 290898 509770 291134
rect 510006 290898 540490 291134
rect 540726 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 33610 273454
rect 33846 273218 64330 273454
rect 64566 273218 95050 273454
rect 95286 273218 125770 273454
rect 126006 273218 156490 273454
rect 156726 273218 187210 273454
rect 187446 273218 217930 273454
rect 218166 273218 248650 273454
rect 248886 273218 279370 273454
rect 279606 273218 310090 273454
rect 310326 273218 340810 273454
rect 341046 273218 371530 273454
rect 371766 273218 402250 273454
rect 402486 273218 432970 273454
rect 433206 273218 463690 273454
rect 463926 273218 494410 273454
rect 494646 273218 525130 273454
rect 525366 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 33610 273134
rect 33846 272898 64330 273134
rect 64566 272898 95050 273134
rect 95286 272898 125770 273134
rect 126006 272898 156490 273134
rect 156726 272898 187210 273134
rect 187446 272898 217930 273134
rect 218166 272898 248650 273134
rect 248886 272898 279370 273134
rect 279606 272898 310090 273134
rect 310326 272898 340810 273134
rect 341046 272898 371530 273134
rect 371766 272898 402250 273134
rect 402486 272898 432970 273134
rect 433206 272898 463690 273134
rect 463926 272898 494410 273134
rect 494646 272898 525130 273134
rect 525366 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 18250 255454
rect 18486 255218 48970 255454
rect 49206 255218 79690 255454
rect 79926 255218 110410 255454
rect 110646 255218 141130 255454
rect 141366 255218 171850 255454
rect 172086 255218 202570 255454
rect 202806 255218 233290 255454
rect 233526 255218 264010 255454
rect 264246 255218 294730 255454
rect 294966 255218 325450 255454
rect 325686 255218 356170 255454
rect 356406 255218 386890 255454
rect 387126 255218 417610 255454
rect 417846 255218 448330 255454
rect 448566 255218 479050 255454
rect 479286 255218 509770 255454
rect 510006 255218 540490 255454
rect 540726 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 18250 255134
rect 18486 254898 48970 255134
rect 49206 254898 79690 255134
rect 79926 254898 110410 255134
rect 110646 254898 141130 255134
rect 141366 254898 171850 255134
rect 172086 254898 202570 255134
rect 202806 254898 233290 255134
rect 233526 254898 264010 255134
rect 264246 254898 294730 255134
rect 294966 254898 325450 255134
rect 325686 254898 356170 255134
rect 356406 254898 386890 255134
rect 387126 254898 417610 255134
rect 417846 254898 448330 255134
rect 448566 254898 479050 255134
rect 479286 254898 509770 255134
rect 510006 254898 540490 255134
rect 540726 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 33610 237454
rect 33846 237218 64330 237454
rect 64566 237218 95050 237454
rect 95286 237218 125770 237454
rect 126006 237218 156490 237454
rect 156726 237218 187210 237454
rect 187446 237218 217930 237454
rect 218166 237218 248650 237454
rect 248886 237218 279370 237454
rect 279606 237218 310090 237454
rect 310326 237218 340810 237454
rect 341046 237218 371530 237454
rect 371766 237218 402250 237454
rect 402486 237218 432970 237454
rect 433206 237218 463690 237454
rect 463926 237218 494410 237454
rect 494646 237218 525130 237454
rect 525366 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 33610 237134
rect 33846 236898 64330 237134
rect 64566 236898 95050 237134
rect 95286 236898 125770 237134
rect 126006 236898 156490 237134
rect 156726 236898 187210 237134
rect 187446 236898 217930 237134
rect 218166 236898 248650 237134
rect 248886 236898 279370 237134
rect 279606 236898 310090 237134
rect 310326 236898 340810 237134
rect 341046 236898 371530 237134
rect 371766 236898 402250 237134
rect 402486 236898 432970 237134
rect 433206 236898 463690 237134
rect 463926 236898 494410 237134
rect 494646 236898 525130 237134
rect 525366 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 18250 219454
rect 18486 219218 48970 219454
rect 49206 219218 79690 219454
rect 79926 219218 110410 219454
rect 110646 219218 141130 219454
rect 141366 219218 171850 219454
rect 172086 219218 202570 219454
rect 202806 219218 233290 219454
rect 233526 219218 264010 219454
rect 264246 219218 294730 219454
rect 294966 219218 325450 219454
rect 325686 219218 356170 219454
rect 356406 219218 386890 219454
rect 387126 219218 417610 219454
rect 417846 219218 448330 219454
rect 448566 219218 479050 219454
rect 479286 219218 509770 219454
rect 510006 219218 540490 219454
rect 540726 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 18250 219134
rect 18486 218898 48970 219134
rect 49206 218898 79690 219134
rect 79926 218898 110410 219134
rect 110646 218898 141130 219134
rect 141366 218898 171850 219134
rect 172086 218898 202570 219134
rect 202806 218898 233290 219134
rect 233526 218898 264010 219134
rect 264246 218898 294730 219134
rect 294966 218898 325450 219134
rect 325686 218898 356170 219134
rect 356406 218898 386890 219134
rect 387126 218898 417610 219134
rect 417846 218898 448330 219134
rect 448566 218898 479050 219134
rect 479286 218898 509770 219134
rect 510006 218898 540490 219134
rect 540726 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 33610 201454
rect 33846 201218 64330 201454
rect 64566 201218 95050 201454
rect 95286 201218 125770 201454
rect 126006 201218 156490 201454
rect 156726 201218 187210 201454
rect 187446 201218 217930 201454
rect 218166 201218 248650 201454
rect 248886 201218 279370 201454
rect 279606 201218 310090 201454
rect 310326 201218 340810 201454
rect 341046 201218 371530 201454
rect 371766 201218 402250 201454
rect 402486 201218 432970 201454
rect 433206 201218 463690 201454
rect 463926 201218 494410 201454
rect 494646 201218 525130 201454
rect 525366 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 33610 201134
rect 33846 200898 64330 201134
rect 64566 200898 95050 201134
rect 95286 200898 125770 201134
rect 126006 200898 156490 201134
rect 156726 200898 187210 201134
rect 187446 200898 217930 201134
rect 218166 200898 248650 201134
rect 248886 200898 279370 201134
rect 279606 200898 310090 201134
rect 310326 200898 340810 201134
rect 341046 200898 371530 201134
rect 371766 200898 402250 201134
rect 402486 200898 432970 201134
rect 433206 200898 463690 201134
rect 463926 200898 494410 201134
rect 494646 200898 525130 201134
rect 525366 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 18250 183454
rect 18486 183218 48970 183454
rect 49206 183218 79690 183454
rect 79926 183218 110410 183454
rect 110646 183218 141130 183454
rect 141366 183218 171850 183454
rect 172086 183218 202570 183454
rect 202806 183218 233290 183454
rect 233526 183218 264010 183454
rect 264246 183218 294730 183454
rect 294966 183218 325450 183454
rect 325686 183218 356170 183454
rect 356406 183218 386890 183454
rect 387126 183218 417610 183454
rect 417846 183218 448330 183454
rect 448566 183218 479050 183454
rect 479286 183218 509770 183454
rect 510006 183218 540490 183454
rect 540726 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 18250 183134
rect 18486 182898 48970 183134
rect 49206 182898 79690 183134
rect 79926 182898 110410 183134
rect 110646 182898 141130 183134
rect 141366 182898 171850 183134
rect 172086 182898 202570 183134
rect 202806 182898 233290 183134
rect 233526 182898 264010 183134
rect 264246 182898 294730 183134
rect 294966 182898 325450 183134
rect 325686 182898 356170 183134
rect 356406 182898 386890 183134
rect 387126 182898 417610 183134
rect 417846 182898 448330 183134
rect 448566 182898 479050 183134
rect 479286 182898 509770 183134
rect 510006 182898 540490 183134
rect 540726 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 33610 165454
rect 33846 165218 64330 165454
rect 64566 165218 95050 165454
rect 95286 165218 125770 165454
rect 126006 165218 156490 165454
rect 156726 165218 187210 165454
rect 187446 165218 217930 165454
rect 218166 165218 248650 165454
rect 248886 165218 279370 165454
rect 279606 165218 310090 165454
rect 310326 165218 340810 165454
rect 341046 165218 371530 165454
rect 371766 165218 402250 165454
rect 402486 165218 432970 165454
rect 433206 165218 463690 165454
rect 463926 165218 494410 165454
rect 494646 165218 525130 165454
rect 525366 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 33610 165134
rect 33846 164898 64330 165134
rect 64566 164898 95050 165134
rect 95286 164898 125770 165134
rect 126006 164898 156490 165134
rect 156726 164898 187210 165134
rect 187446 164898 217930 165134
rect 218166 164898 248650 165134
rect 248886 164898 279370 165134
rect 279606 164898 310090 165134
rect 310326 164898 340810 165134
rect 341046 164898 371530 165134
rect 371766 164898 402250 165134
rect 402486 164898 432970 165134
rect 433206 164898 463690 165134
rect 463926 164898 494410 165134
rect 494646 164898 525130 165134
rect 525366 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 18250 147454
rect 18486 147218 48970 147454
rect 49206 147218 79690 147454
rect 79926 147218 110410 147454
rect 110646 147218 141130 147454
rect 141366 147218 171850 147454
rect 172086 147218 202570 147454
rect 202806 147218 233290 147454
rect 233526 147218 264010 147454
rect 264246 147218 294730 147454
rect 294966 147218 325450 147454
rect 325686 147218 356170 147454
rect 356406 147218 386890 147454
rect 387126 147218 417610 147454
rect 417846 147218 448330 147454
rect 448566 147218 479050 147454
rect 479286 147218 509770 147454
rect 510006 147218 540490 147454
rect 540726 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 18250 147134
rect 18486 146898 48970 147134
rect 49206 146898 79690 147134
rect 79926 146898 110410 147134
rect 110646 146898 141130 147134
rect 141366 146898 171850 147134
rect 172086 146898 202570 147134
rect 202806 146898 233290 147134
rect 233526 146898 264010 147134
rect 264246 146898 294730 147134
rect 294966 146898 325450 147134
rect 325686 146898 356170 147134
rect 356406 146898 386890 147134
rect 387126 146898 417610 147134
rect 417846 146898 448330 147134
rect 448566 146898 479050 147134
rect 479286 146898 509770 147134
rect 510006 146898 540490 147134
rect 540726 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 33610 129454
rect 33846 129218 64330 129454
rect 64566 129218 95050 129454
rect 95286 129218 125770 129454
rect 126006 129218 156490 129454
rect 156726 129218 187210 129454
rect 187446 129218 217930 129454
rect 218166 129218 248650 129454
rect 248886 129218 279370 129454
rect 279606 129218 310090 129454
rect 310326 129218 340810 129454
rect 341046 129218 371530 129454
rect 371766 129218 402250 129454
rect 402486 129218 432970 129454
rect 433206 129218 463690 129454
rect 463926 129218 494410 129454
rect 494646 129218 525130 129454
rect 525366 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 33610 129134
rect 33846 128898 64330 129134
rect 64566 128898 95050 129134
rect 95286 128898 125770 129134
rect 126006 128898 156490 129134
rect 156726 128898 187210 129134
rect 187446 128898 217930 129134
rect 218166 128898 248650 129134
rect 248886 128898 279370 129134
rect 279606 128898 310090 129134
rect 310326 128898 340810 129134
rect 341046 128898 371530 129134
rect 371766 128898 402250 129134
rect 402486 128898 432970 129134
rect 433206 128898 463690 129134
rect 463926 128898 494410 129134
rect 494646 128898 525130 129134
rect 525366 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 18250 111454
rect 18486 111218 48970 111454
rect 49206 111218 79690 111454
rect 79926 111218 110410 111454
rect 110646 111218 141130 111454
rect 141366 111218 171850 111454
rect 172086 111218 202570 111454
rect 202806 111218 233290 111454
rect 233526 111218 264010 111454
rect 264246 111218 294730 111454
rect 294966 111218 325450 111454
rect 325686 111218 356170 111454
rect 356406 111218 386890 111454
rect 387126 111218 417610 111454
rect 417846 111218 448330 111454
rect 448566 111218 479050 111454
rect 479286 111218 509770 111454
rect 510006 111218 540490 111454
rect 540726 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 18250 111134
rect 18486 110898 48970 111134
rect 49206 110898 79690 111134
rect 79926 110898 110410 111134
rect 110646 110898 141130 111134
rect 141366 110898 171850 111134
rect 172086 110898 202570 111134
rect 202806 110898 233290 111134
rect 233526 110898 264010 111134
rect 264246 110898 294730 111134
rect 294966 110898 325450 111134
rect 325686 110898 356170 111134
rect 356406 110898 386890 111134
rect 387126 110898 417610 111134
rect 417846 110898 448330 111134
rect 448566 110898 479050 111134
rect 479286 110898 509770 111134
rect 510006 110898 540490 111134
rect 540726 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 33610 93454
rect 33846 93218 64330 93454
rect 64566 93218 95050 93454
rect 95286 93218 125770 93454
rect 126006 93218 156490 93454
rect 156726 93218 187210 93454
rect 187446 93218 217930 93454
rect 218166 93218 248650 93454
rect 248886 93218 279370 93454
rect 279606 93218 310090 93454
rect 310326 93218 340810 93454
rect 341046 93218 371530 93454
rect 371766 93218 402250 93454
rect 402486 93218 432970 93454
rect 433206 93218 463690 93454
rect 463926 93218 494410 93454
rect 494646 93218 525130 93454
rect 525366 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 33610 93134
rect 33846 92898 64330 93134
rect 64566 92898 95050 93134
rect 95286 92898 125770 93134
rect 126006 92898 156490 93134
rect 156726 92898 187210 93134
rect 187446 92898 217930 93134
rect 218166 92898 248650 93134
rect 248886 92898 279370 93134
rect 279606 92898 310090 93134
rect 310326 92898 340810 93134
rect 341046 92898 371530 93134
rect 371766 92898 402250 93134
rect 402486 92898 432970 93134
rect 433206 92898 463690 93134
rect 463926 92898 494410 93134
rect 494646 92898 525130 93134
rect 525366 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 18250 75454
rect 18486 75218 48970 75454
rect 49206 75218 79690 75454
rect 79926 75218 110410 75454
rect 110646 75218 141130 75454
rect 141366 75218 171850 75454
rect 172086 75218 202570 75454
rect 202806 75218 233290 75454
rect 233526 75218 264010 75454
rect 264246 75218 294730 75454
rect 294966 75218 325450 75454
rect 325686 75218 356170 75454
rect 356406 75218 386890 75454
rect 387126 75218 417610 75454
rect 417846 75218 448330 75454
rect 448566 75218 479050 75454
rect 479286 75218 509770 75454
rect 510006 75218 540490 75454
rect 540726 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 18250 75134
rect 18486 74898 48970 75134
rect 49206 74898 79690 75134
rect 79926 74898 110410 75134
rect 110646 74898 141130 75134
rect 141366 74898 171850 75134
rect 172086 74898 202570 75134
rect 202806 74898 233290 75134
rect 233526 74898 264010 75134
rect 264246 74898 294730 75134
rect 294966 74898 325450 75134
rect 325686 74898 356170 75134
rect 356406 74898 386890 75134
rect 387126 74898 417610 75134
rect 417846 74898 448330 75134
rect 448566 74898 479050 75134
rect 479286 74898 509770 75134
rect 510006 74898 540490 75134
rect 540726 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 33610 57454
rect 33846 57218 64330 57454
rect 64566 57218 95050 57454
rect 95286 57218 125770 57454
rect 126006 57218 156490 57454
rect 156726 57218 187210 57454
rect 187446 57218 217930 57454
rect 218166 57218 248650 57454
rect 248886 57218 279370 57454
rect 279606 57218 310090 57454
rect 310326 57218 340810 57454
rect 341046 57218 371530 57454
rect 371766 57218 402250 57454
rect 402486 57218 432970 57454
rect 433206 57218 463690 57454
rect 463926 57218 494410 57454
rect 494646 57218 525130 57454
rect 525366 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 33610 57134
rect 33846 56898 64330 57134
rect 64566 56898 95050 57134
rect 95286 56898 125770 57134
rect 126006 56898 156490 57134
rect 156726 56898 187210 57134
rect 187446 56898 217930 57134
rect 218166 56898 248650 57134
rect 248886 56898 279370 57134
rect 279606 56898 310090 57134
rect 310326 56898 340810 57134
rect 341046 56898 371530 57134
rect 371766 56898 402250 57134
rect 402486 56898 432970 57134
rect 433206 56898 463690 57134
rect 463926 56898 494410 57134
rect 494646 56898 525130 57134
rect 525366 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 14000 0 1 50000
box 13 0 540000 620000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 48000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 672000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 672000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 672000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 672000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 672000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 672000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 672000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 672000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 672000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 672000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 672000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 672000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 672000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 672000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 672000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 48000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 672000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 672000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 672000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 672000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 672000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 672000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 672000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 672000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 672000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 672000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 672000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 672000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 672000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 672000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 672000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 48000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 672000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 672000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 672000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 672000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 672000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 672000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 672000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 672000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 672000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 672000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 672000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 672000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 672000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 672000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 672000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 48000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 672000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 672000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 672000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 672000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 672000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 672000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 672000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 672000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 672000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 672000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 672000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 672000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 672000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 672000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 672000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 672000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 48000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 672000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 672000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 672000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 672000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 672000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 672000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 672000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 672000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 672000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 672000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 672000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 672000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 672000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 672000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 672000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 48000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 672000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 672000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 672000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 672000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 672000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 672000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 672000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 672000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 672000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 672000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 672000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 672000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 672000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 672000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 672000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 48000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 672000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 672000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 672000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 672000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 672000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 672000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 672000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 672000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 672000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 672000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 672000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 672000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 672000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 672000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 672000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 48000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 672000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 672000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 672000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 672000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 672000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 672000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 672000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 672000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 672000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 672000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 672000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 672000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 672000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 672000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 672000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
