magic
tech sky130A
magscale 1 2
timestamp 1650987940
<< obsli1 >>
rect 1104 2159 538844 617457
<< obsm1 >>
rect 1104 1980 539474 617488
<< metal2 >>
rect 2318 619200 2374 620000
rect 7010 619200 7066 620000
rect 11702 619200 11758 620000
rect 16394 619200 16450 620000
rect 21086 619200 21142 620000
rect 25778 619200 25834 620000
rect 30470 619200 30526 620000
rect 35162 619200 35218 620000
rect 39854 619200 39910 620000
rect 44546 619200 44602 620000
rect 49238 619200 49294 620000
rect 53930 619200 53986 620000
rect 58622 619200 58678 620000
rect 63314 619200 63370 620000
rect 68006 619200 68062 620000
rect 72698 619200 72754 620000
rect 77390 619200 77446 620000
rect 82082 619200 82138 620000
rect 86774 619200 86830 620000
rect 91466 619200 91522 620000
rect 96158 619200 96214 620000
rect 100850 619200 100906 620000
rect 105542 619200 105598 620000
rect 110326 619200 110382 620000
rect 115018 619200 115074 620000
rect 119710 619200 119766 620000
rect 124402 619200 124458 620000
rect 129094 619200 129150 620000
rect 133786 619200 133842 620000
rect 138478 619200 138534 620000
rect 143170 619200 143226 620000
rect 147862 619200 147918 620000
rect 152554 619200 152610 620000
rect 157246 619200 157302 620000
rect 161938 619200 161994 620000
rect 166630 619200 166686 620000
rect 171322 619200 171378 620000
rect 176014 619200 176070 620000
rect 180706 619200 180762 620000
rect 185398 619200 185454 620000
rect 190090 619200 190146 620000
rect 194782 619200 194838 620000
rect 199474 619200 199530 620000
rect 204166 619200 204222 620000
rect 208858 619200 208914 620000
rect 213550 619200 213606 620000
rect 218334 619200 218390 620000
rect 223026 619200 223082 620000
rect 227718 619200 227774 620000
rect 232410 619200 232466 620000
rect 237102 619200 237158 620000
rect 241794 619200 241850 620000
rect 246486 619200 246542 620000
rect 251178 619200 251234 620000
rect 255870 619200 255926 620000
rect 260562 619200 260618 620000
rect 265254 619200 265310 620000
rect 269946 619200 270002 620000
rect 274638 619200 274694 620000
rect 279330 619200 279386 620000
rect 284022 619200 284078 620000
rect 288714 619200 288770 620000
rect 293406 619200 293462 620000
rect 298098 619200 298154 620000
rect 302790 619200 302846 620000
rect 307482 619200 307538 620000
rect 312174 619200 312230 620000
rect 316866 619200 316922 620000
rect 321558 619200 321614 620000
rect 326342 619200 326398 620000
rect 331034 619200 331090 620000
rect 335726 619200 335782 620000
rect 340418 619200 340474 620000
rect 345110 619200 345166 620000
rect 349802 619200 349858 620000
rect 354494 619200 354550 620000
rect 359186 619200 359242 620000
rect 363878 619200 363934 620000
rect 368570 619200 368626 620000
rect 373262 619200 373318 620000
rect 377954 619200 378010 620000
rect 382646 619200 382702 620000
rect 387338 619200 387394 620000
rect 392030 619200 392086 620000
rect 396722 619200 396778 620000
rect 401414 619200 401470 620000
rect 406106 619200 406162 620000
rect 410798 619200 410854 620000
rect 415490 619200 415546 620000
rect 420182 619200 420238 620000
rect 424874 619200 424930 620000
rect 429566 619200 429622 620000
rect 434350 619200 434406 620000
rect 439042 619200 439098 620000
rect 443734 619200 443790 620000
rect 448426 619200 448482 620000
rect 453118 619200 453174 620000
rect 457810 619200 457866 620000
rect 462502 619200 462558 620000
rect 467194 619200 467250 620000
rect 471886 619200 471942 620000
rect 476578 619200 476634 620000
rect 481270 619200 481326 620000
rect 485962 619200 486018 620000
rect 490654 619200 490710 620000
rect 495346 619200 495402 620000
rect 500038 619200 500094 620000
rect 504730 619200 504786 620000
rect 509422 619200 509478 620000
rect 514114 619200 514170 620000
rect 518806 619200 518862 620000
rect 523498 619200 523554 620000
rect 528190 619200 528246 620000
rect 532882 619200 532938 620000
rect 537574 619200 537630 620000
rect 478 0 534 800
rect 1490 0 1546 800
rect 2594 0 2650 800
rect 3698 0 3754 800
rect 4802 0 4858 800
rect 5906 0 5962 800
rect 7010 0 7066 800
rect 8114 0 8170 800
rect 9218 0 9274 800
rect 10322 0 10378 800
rect 11426 0 11482 800
rect 12438 0 12494 800
rect 13542 0 13598 800
rect 14646 0 14702 800
rect 15750 0 15806 800
rect 16854 0 16910 800
rect 17958 0 18014 800
rect 19062 0 19118 800
rect 20166 0 20222 800
rect 21270 0 21326 800
rect 22374 0 22430 800
rect 23478 0 23534 800
rect 24490 0 24546 800
rect 25594 0 25650 800
rect 26698 0 26754 800
rect 27802 0 27858 800
rect 28906 0 28962 800
rect 30010 0 30066 800
rect 31114 0 31170 800
rect 32218 0 32274 800
rect 33322 0 33378 800
rect 34426 0 34482 800
rect 35530 0 35586 800
rect 36542 0 36598 800
rect 37646 0 37702 800
rect 38750 0 38806 800
rect 39854 0 39910 800
rect 40958 0 41014 800
rect 42062 0 42118 800
rect 43166 0 43222 800
rect 44270 0 44326 800
rect 45374 0 45430 800
rect 46478 0 46534 800
rect 47490 0 47546 800
rect 48594 0 48650 800
rect 49698 0 49754 800
rect 50802 0 50858 800
rect 51906 0 51962 800
rect 53010 0 53066 800
rect 54114 0 54170 800
rect 55218 0 55274 800
rect 56322 0 56378 800
rect 57426 0 57482 800
rect 58530 0 58586 800
rect 59542 0 59598 800
rect 60646 0 60702 800
rect 61750 0 61806 800
rect 62854 0 62910 800
rect 63958 0 64014 800
rect 65062 0 65118 800
rect 66166 0 66222 800
rect 67270 0 67326 800
rect 68374 0 68430 800
rect 69478 0 69534 800
rect 70582 0 70638 800
rect 71594 0 71650 800
rect 72698 0 72754 800
rect 73802 0 73858 800
rect 74906 0 74962 800
rect 76010 0 76066 800
rect 77114 0 77170 800
rect 78218 0 78274 800
rect 79322 0 79378 800
rect 80426 0 80482 800
rect 81530 0 81586 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84750 0 84806 800
rect 85854 0 85910 800
rect 86958 0 87014 800
rect 88062 0 88118 800
rect 89166 0 89222 800
rect 90270 0 90326 800
rect 91374 0 91430 800
rect 92478 0 92534 800
rect 93582 0 93638 800
rect 94594 0 94650 800
rect 95698 0 95754 800
rect 96802 0 96858 800
rect 97906 0 97962 800
rect 99010 0 99066 800
rect 100114 0 100170 800
rect 101218 0 101274 800
rect 102322 0 102378 800
rect 103426 0 103482 800
rect 104530 0 104586 800
rect 105634 0 105690 800
rect 106646 0 106702 800
rect 107750 0 107806 800
rect 108854 0 108910 800
rect 109958 0 110014 800
rect 111062 0 111118 800
rect 112166 0 112222 800
rect 113270 0 113326 800
rect 114374 0 114430 800
rect 115478 0 115534 800
rect 116582 0 116638 800
rect 117686 0 117742 800
rect 118698 0 118754 800
rect 119802 0 119858 800
rect 120906 0 120962 800
rect 122010 0 122066 800
rect 123114 0 123170 800
rect 124218 0 124274 800
rect 125322 0 125378 800
rect 126426 0 126482 800
rect 127530 0 127586 800
rect 128634 0 128690 800
rect 129646 0 129702 800
rect 130750 0 130806 800
rect 131854 0 131910 800
rect 132958 0 133014 800
rect 134062 0 134118 800
rect 135166 0 135222 800
rect 136270 0 136326 800
rect 137374 0 137430 800
rect 138478 0 138534 800
rect 139582 0 139638 800
rect 140686 0 140742 800
rect 141698 0 141754 800
rect 142802 0 142858 800
rect 143906 0 143962 800
rect 145010 0 145066 800
rect 146114 0 146170 800
rect 147218 0 147274 800
rect 148322 0 148378 800
rect 149426 0 149482 800
rect 150530 0 150586 800
rect 151634 0 151690 800
rect 152738 0 152794 800
rect 153750 0 153806 800
rect 154854 0 154910 800
rect 155958 0 156014 800
rect 157062 0 157118 800
rect 158166 0 158222 800
rect 159270 0 159326 800
rect 160374 0 160430 800
rect 161478 0 161534 800
rect 162582 0 162638 800
rect 163686 0 163742 800
rect 164790 0 164846 800
rect 165802 0 165858 800
rect 166906 0 166962 800
rect 168010 0 168066 800
rect 169114 0 169170 800
rect 170218 0 170274 800
rect 171322 0 171378 800
rect 172426 0 172482 800
rect 173530 0 173586 800
rect 174634 0 174690 800
rect 175738 0 175794 800
rect 176750 0 176806 800
rect 177854 0 177910 800
rect 178958 0 179014 800
rect 180062 0 180118 800
rect 181166 0 181222 800
rect 182270 0 182326 800
rect 183374 0 183430 800
rect 184478 0 184534 800
rect 185582 0 185638 800
rect 186686 0 186742 800
rect 187790 0 187846 800
rect 188802 0 188858 800
rect 189906 0 189962 800
rect 191010 0 191066 800
rect 192114 0 192170 800
rect 193218 0 193274 800
rect 194322 0 194378 800
rect 195426 0 195482 800
rect 196530 0 196586 800
rect 197634 0 197690 800
rect 198738 0 198794 800
rect 199842 0 199898 800
rect 200854 0 200910 800
rect 201958 0 202014 800
rect 203062 0 203118 800
rect 204166 0 204222 800
rect 205270 0 205326 800
rect 206374 0 206430 800
rect 207478 0 207534 800
rect 208582 0 208638 800
rect 209686 0 209742 800
rect 210790 0 210846 800
rect 211802 0 211858 800
rect 212906 0 212962 800
rect 214010 0 214066 800
rect 215114 0 215170 800
rect 216218 0 216274 800
rect 217322 0 217378 800
rect 218426 0 218482 800
rect 219530 0 219586 800
rect 220634 0 220690 800
rect 221738 0 221794 800
rect 222842 0 222898 800
rect 223854 0 223910 800
rect 224958 0 225014 800
rect 226062 0 226118 800
rect 227166 0 227222 800
rect 228270 0 228326 800
rect 229374 0 229430 800
rect 230478 0 230534 800
rect 231582 0 231638 800
rect 232686 0 232742 800
rect 233790 0 233846 800
rect 234894 0 234950 800
rect 235906 0 235962 800
rect 237010 0 237066 800
rect 238114 0 238170 800
rect 239218 0 239274 800
rect 240322 0 240378 800
rect 241426 0 241482 800
rect 242530 0 242586 800
rect 243634 0 243690 800
rect 244738 0 244794 800
rect 245842 0 245898 800
rect 246946 0 247002 800
rect 247958 0 248014 800
rect 249062 0 249118 800
rect 250166 0 250222 800
rect 251270 0 251326 800
rect 252374 0 252430 800
rect 253478 0 253534 800
rect 254582 0 254638 800
rect 255686 0 255742 800
rect 256790 0 256846 800
rect 257894 0 257950 800
rect 258906 0 258962 800
rect 260010 0 260066 800
rect 261114 0 261170 800
rect 262218 0 262274 800
rect 263322 0 263378 800
rect 264426 0 264482 800
rect 265530 0 265586 800
rect 266634 0 266690 800
rect 267738 0 267794 800
rect 268842 0 268898 800
rect 269946 0 270002 800
rect 270958 0 271014 800
rect 272062 0 272118 800
rect 273166 0 273222 800
rect 274270 0 274326 800
rect 275374 0 275430 800
rect 276478 0 276534 800
rect 277582 0 277638 800
rect 278686 0 278742 800
rect 279790 0 279846 800
rect 280894 0 280950 800
rect 281998 0 282054 800
rect 283010 0 283066 800
rect 284114 0 284170 800
rect 285218 0 285274 800
rect 286322 0 286378 800
rect 287426 0 287482 800
rect 288530 0 288586 800
rect 289634 0 289690 800
rect 290738 0 290794 800
rect 291842 0 291898 800
rect 292946 0 293002 800
rect 293958 0 294014 800
rect 295062 0 295118 800
rect 296166 0 296222 800
rect 297270 0 297326 800
rect 298374 0 298430 800
rect 299478 0 299534 800
rect 300582 0 300638 800
rect 301686 0 301742 800
rect 302790 0 302846 800
rect 303894 0 303950 800
rect 304998 0 305054 800
rect 306010 0 306066 800
rect 307114 0 307170 800
rect 308218 0 308274 800
rect 309322 0 309378 800
rect 310426 0 310482 800
rect 311530 0 311586 800
rect 312634 0 312690 800
rect 313738 0 313794 800
rect 314842 0 314898 800
rect 315946 0 316002 800
rect 317050 0 317106 800
rect 318062 0 318118 800
rect 319166 0 319222 800
rect 320270 0 320326 800
rect 321374 0 321430 800
rect 322478 0 322534 800
rect 323582 0 323638 800
rect 324686 0 324742 800
rect 325790 0 325846 800
rect 326894 0 326950 800
rect 327998 0 328054 800
rect 329102 0 329158 800
rect 330114 0 330170 800
rect 331218 0 331274 800
rect 332322 0 332378 800
rect 333426 0 333482 800
rect 334530 0 334586 800
rect 335634 0 335690 800
rect 336738 0 336794 800
rect 337842 0 337898 800
rect 338946 0 339002 800
rect 340050 0 340106 800
rect 341062 0 341118 800
rect 342166 0 342222 800
rect 343270 0 343326 800
rect 344374 0 344430 800
rect 345478 0 345534 800
rect 346582 0 346638 800
rect 347686 0 347742 800
rect 348790 0 348846 800
rect 349894 0 349950 800
rect 350998 0 351054 800
rect 352102 0 352158 800
rect 353114 0 353170 800
rect 354218 0 354274 800
rect 355322 0 355378 800
rect 356426 0 356482 800
rect 357530 0 357586 800
rect 358634 0 358690 800
rect 359738 0 359794 800
rect 360842 0 360898 800
rect 361946 0 362002 800
rect 363050 0 363106 800
rect 364154 0 364210 800
rect 365166 0 365222 800
rect 366270 0 366326 800
rect 367374 0 367430 800
rect 368478 0 368534 800
rect 369582 0 369638 800
rect 370686 0 370742 800
rect 371790 0 371846 800
rect 372894 0 372950 800
rect 373998 0 374054 800
rect 375102 0 375158 800
rect 376114 0 376170 800
rect 377218 0 377274 800
rect 378322 0 378378 800
rect 379426 0 379482 800
rect 380530 0 380586 800
rect 381634 0 381690 800
rect 382738 0 382794 800
rect 383842 0 383898 800
rect 384946 0 385002 800
rect 386050 0 386106 800
rect 387154 0 387210 800
rect 388166 0 388222 800
rect 389270 0 389326 800
rect 390374 0 390430 800
rect 391478 0 391534 800
rect 392582 0 392638 800
rect 393686 0 393742 800
rect 394790 0 394846 800
rect 395894 0 395950 800
rect 396998 0 397054 800
rect 398102 0 398158 800
rect 399206 0 399262 800
rect 400218 0 400274 800
rect 401322 0 401378 800
rect 402426 0 402482 800
rect 403530 0 403586 800
rect 404634 0 404690 800
rect 405738 0 405794 800
rect 406842 0 406898 800
rect 407946 0 408002 800
rect 409050 0 409106 800
rect 410154 0 410210 800
rect 411258 0 411314 800
rect 412270 0 412326 800
rect 413374 0 413430 800
rect 414478 0 414534 800
rect 415582 0 415638 800
rect 416686 0 416742 800
rect 417790 0 417846 800
rect 418894 0 418950 800
rect 419998 0 420054 800
rect 421102 0 421158 800
rect 422206 0 422262 800
rect 423218 0 423274 800
rect 424322 0 424378 800
rect 425426 0 425482 800
rect 426530 0 426586 800
rect 427634 0 427690 800
rect 428738 0 428794 800
rect 429842 0 429898 800
rect 430946 0 431002 800
rect 432050 0 432106 800
rect 433154 0 433210 800
rect 434258 0 434314 800
rect 435270 0 435326 800
rect 436374 0 436430 800
rect 437478 0 437534 800
rect 438582 0 438638 800
rect 439686 0 439742 800
rect 440790 0 440846 800
rect 441894 0 441950 800
rect 442998 0 443054 800
rect 444102 0 444158 800
rect 445206 0 445262 800
rect 446310 0 446366 800
rect 447322 0 447378 800
rect 448426 0 448482 800
rect 449530 0 449586 800
rect 450634 0 450690 800
rect 451738 0 451794 800
rect 452842 0 452898 800
rect 453946 0 454002 800
rect 455050 0 455106 800
rect 456154 0 456210 800
rect 457258 0 457314 800
rect 458270 0 458326 800
rect 459374 0 459430 800
rect 460478 0 460534 800
rect 461582 0 461638 800
rect 462686 0 462742 800
rect 463790 0 463846 800
rect 464894 0 464950 800
rect 465998 0 466054 800
rect 467102 0 467158 800
rect 468206 0 468262 800
rect 469310 0 469366 800
rect 470322 0 470378 800
rect 471426 0 471482 800
rect 472530 0 472586 800
rect 473634 0 473690 800
rect 474738 0 474794 800
rect 475842 0 475898 800
rect 476946 0 477002 800
rect 478050 0 478106 800
rect 479154 0 479210 800
rect 480258 0 480314 800
rect 481362 0 481418 800
rect 482374 0 482430 800
rect 483478 0 483534 800
rect 484582 0 484638 800
rect 485686 0 485742 800
rect 486790 0 486846 800
rect 487894 0 487950 800
rect 488998 0 489054 800
rect 490102 0 490158 800
rect 491206 0 491262 800
rect 492310 0 492366 800
rect 493414 0 493470 800
rect 494426 0 494482 800
rect 495530 0 495586 800
rect 496634 0 496690 800
rect 497738 0 497794 800
rect 498842 0 498898 800
rect 499946 0 500002 800
rect 501050 0 501106 800
rect 502154 0 502210 800
rect 503258 0 503314 800
rect 504362 0 504418 800
rect 505374 0 505430 800
rect 506478 0 506534 800
rect 507582 0 507638 800
rect 508686 0 508742 800
rect 509790 0 509846 800
rect 510894 0 510950 800
rect 511998 0 512054 800
rect 513102 0 513158 800
rect 514206 0 514262 800
rect 515310 0 515366 800
rect 516414 0 516470 800
rect 517426 0 517482 800
rect 518530 0 518586 800
rect 519634 0 519690 800
rect 520738 0 520794 800
rect 521842 0 521898 800
rect 522946 0 523002 800
rect 524050 0 524106 800
rect 525154 0 525210 800
rect 526258 0 526314 800
rect 527362 0 527418 800
rect 528466 0 528522 800
rect 529478 0 529534 800
rect 530582 0 530638 800
rect 531686 0 531742 800
rect 532790 0 532846 800
rect 533894 0 533950 800
rect 534998 0 535054 800
rect 536102 0 536158 800
rect 537206 0 537262 800
rect 538310 0 538366 800
rect 539414 0 539470 800
<< obsm2 >>
rect 18 619144 2262 619200
rect 2430 619144 6954 619200
rect 7122 619144 11646 619200
rect 11814 619144 16338 619200
rect 16506 619144 21030 619200
rect 21198 619144 25722 619200
rect 25890 619144 30414 619200
rect 30582 619144 35106 619200
rect 35274 619144 39798 619200
rect 39966 619144 44490 619200
rect 44658 619144 49182 619200
rect 49350 619144 53874 619200
rect 54042 619144 58566 619200
rect 58734 619144 63258 619200
rect 63426 619144 67950 619200
rect 68118 619144 72642 619200
rect 72810 619144 77334 619200
rect 77502 619144 82026 619200
rect 82194 619144 86718 619200
rect 86886 619144 91410 619200
rect 91578 619144 96102 619200
rect 96270 619144 100794 619200
rect 100962 619144 105486 619200
rect 105654 619144 110270 619200
rect 110438 619144 114962 619200
rect 115130 619144 119654 619200
rect 119822 619144 124346 619200
rect 124514 619144 129038 619200
rect 129206 619144 133730 619200
rect 133898 619144 138422 619200
rect 138590 619144 143114 619200
rect 143282 619144 147806 619200
rect 147974 619144 152498 619200
rect 152666 619144 157190 619200
rect 157358 619144 161882 619200
rect 162050 619144 166574 619200
rect 166742 619144 171266 619200
rect 171434 619144 175958 619200
rect 176126 619144 180650 619200
rect 180818 619144 185342 619200
rect 185510 619144 190034 619200
rect 190202 619144 194726 619200
rect 194894 619144 199418 619200
rect 199586 619144 204110 619200
rect 204278 619144 208802 619200
rect 208970 619144 213494 619200
rect 213662 619144 218278 619200
rect 218446 619144 222970 619200
rect 223138 619144 227662 619200
rect 227830 619144 232354 619200
rect 232522 619144 237046 619200
rect 237214 619144 241738 619200
rect 241906 619144 246430 619200
rect 246598 619144 251122 619200
rect 251290 619144 255814 619200
rect 255982 619144 260506 619200
rect 260674 619144 265198 619200
rect 265366 619144 269890 619200
rect 270058 619144 274582 619200
rect 274750 619144 279274 619200
rect 279442 619144 283966 619200
rect 284134 619144 288658 619200
rect 288826 619144 293350 619200
rect 293518 619144 298042 619200
rect 298210 619144 302734 619200
rect 302902 619144 307426 619200
rect 307594 619144 312118 619200
rect 312286 619144 316810 619200
rect 316978 619144 321502 619200
rect 321670 619144 326286 619200
rect 326454 619144 330978 619200
rect 331146 619144 335670 619200
rect 335838 619144 340362 619200
rect 340530 619144 345054 619200
rect 345222 619144 349746 619200
rect 349914 619144 354438 619200
rect 354606 619144 359130 619200
rect 359298 619144 363822 619200
rect 363990 619144 368514 619200
rect 368682 619144 373206 619200
rect 373374 619144 377898 619200
rect 378066 619144 382590 619200
rect 382758 619144 387282 619200
rect 387450 619144 391974 619200
rect 392142 619144 396666 619200
rect 396834 619144 401358 619200
rect 401526 619144 406050 619200
rect 406218 619144 410742 619200
rect 410910 619144 415434 619200
rect 415602 619144 420126 619200
rect 420294 619144 424818 619200
rect 424986 619144 429510 619200
rect 429678 619144 434294 619200
rect 434462 619144 438986 619200
rect 439154 619144 443678 619200
rect 443846 619144 448370 619200
rect 448538 619144 453062 619200
rect 453230 619144 457754 619200
rect 457922 619144 462446 619200
rect 462614 619144 467138 619200
rect 467306 619144 471830 619200
rect 471998 619144 476522 619200
rect 476690 619144 481214 619200
rect 481382 619144 485906 619200
rect 486074 619144 490598 619200
rect 490766 619144 495290 619200
rect 495458 619144 499982 619200
rect 500150 619144 504674 619200
rect 504842 619144 509366 619200
rect 509534 619144 514058 619200
rect 514226 619144 518750 619200
rect 518918 619144 523442 619200
rect 523610 619144 528134 619200
rect 528302 619144 532826 619200
rect 532994 619144 537518 619200
rect 537686 619144 539468 619200
rect 18 856 539468 619144
rect 18 734 422 856
rect 590 734 1434 856
rect 1602 734 2538 856
rect 2706 734 3642 856
rect 3810 734 4746 856
rect 4914 734 5850 856
rect 6018 734 6954 856
rect 7122 734 8058 856
rect 8226 734 9162 856
rect 9330 734 10266 856
rect 10434 734 11370 856
rect 11538 734 12382 856
rect 12550 734 13486 856
rect 13654 734 14590 856
rect 14758 734 15694 856
rect 15862 734 16798 856
rect 16966 734 17902 856
rect 18070 734 19006 856
rect 19174 734 20110 856
rect 20278 734 21214 856
rect 21382 734 22318 856
rect 22486 734 23422 856
rect 23590 734 24434 856
rect 24602 734 25538 856
rect 25706 734 26642 856
rect 26810 734 27746 856
rect 27914 734 28850 856
rect 29018 734 29954 856
rect 30122 734 31058 856
rect 31226 734 32162 856
rect 32330 734 33266 856
rect 33434 734 34370 856
rect 34538 734 35474 856
rect 35642 734 36486 856
rect 36654 734 37590 856
rect 37758 734 38694 856
rect 38862 734 39798 856
rect 39966 734 40902 856
rect 41070 734 42006 856
rect 42174 734 43110 856
rect 43278 734 44214 856
rect 44382 734 45318 856
rect 45486 734 46422 856
rect 46590 734 47434 856
rect 47602 734 48538 856
rect 48706 734 49642 856
rect 49810 734 50746 856
rect 50914 734 51850 856
rect 52018 734 52954 856
rect 53122 734 54058 856
rect 54226 734 55162 856
rect 55330 734 56266 856
rect 56434 734 57370 856
rect 57538 734 58474 856
rect 58642 734 59486 856
rect 59654 734 60590 856
rect 60758 734 61694 856
rect 61862 734 62798 856
rect 62966 734 63902 856
rect 64070 734 65006 856
rect 65174 734 66110 856
rect 66278 734 67214 856
rect 67382 734 68318 856
rect 68486 734 69422 856
rect 69590 734 70526 856
rect 70694 734 71538 856
rect 71706 734 72642 856
rect 72810 734 73746 856
rect 73914 734 74850 856
rect 75018 734 75954 856
rect 76122 734 77058 856
rect 77226 734 78162 856
rect 78330 734 79266 856
rect 79434 734 80370 856
rect 80538 734 81474 856
rect 81642 734 82578 856
rect 82746 734 83590 856
rect 83758 734 84694 856
rect 84862 734 85798 856
rect 85966 734 86902 856
rect 87070 734 88006 856
rect 88174 734 89110 856
rect 89278 734 90214 856
rect 90382 734 91318 856
rect 91486 734 92422 856
rect 92590 734 93526 856
rect 93694 734 94538 856
rect 94706 734 95642 856
rect 95810 734 96746 856
rect 96914 734 97850 856
rect 98018 734 98954 856
rect 99122 734 100058 856
rect 100226 734 101162 856
rect 101330 734 102266 856
rect 102434 734 103370 856
rect 103538 734 104474 856
rect 104642 734 105578 856
rect 105746 734 106590 856
rect 106758 734 107694 856
rect 107862 734 108798 856
rect 108966 734 109902 856
rect 110070 734 111006 856
rect 111174 734 112110 856
rect 112278 734 113214 856
rect 113382 734 114318 856
rect 114486 734 115422 856
rect 115590 734 116526 856
rect 116694 734 117630 856
rect 117798 734 118642 856
rect 118810 734 119746 856
rect 119914 734 120850 856
rect 121018 734 121954 856
rect 122122 734 123058 856
rect 123226 734 124162 856
rect 124330 734 125266 856
rect 125434 734 126370 856
rect 126538 734 127474 856
rect 127642 734 128578 856
rect 128746 734 129590 856
rect 129758 734 130694 856
rect 130862 734 131798 856
rect 131966 734 132902 856
rect 133070 734 134006 856
rect 134174 734 135110 856
rect 135278 734 136214 856
rect 136382 734 137318 856
rect 137486 734 138422 856
rect 138590 734 139526 856
rect 139694 734 140630 856
rect 140798 734 141642 856
rect 141810 734 142746 856
rect 142914 734 143850 856
rect 144018 734 144954 856
rect 145122 734 146058 856
rect 146226 734 147162 856
rect 147330 734 148266 856
rect 148434 734 149370 856
rect 149538 734 150474 856
rect 150642 734 151578 856
rect 151746 734 152682 856
rect 152850 734 153694 856
rect 153862 734 154798 856
rect 154966 734 155902 856
rect 156070 734 157006 856
rect 157174 734 158110 856
rect 158278 734 159214 856
rect 159382 734 160318 856
rect 160486 734 161422 856
rect 161590 734 162526 856
rect 162694 734 163630 856
rect 163798 734 164734 856
rect 164902 734 165746 856
rect 165914 734 166850 856
rect 167018 734 167954 856
rect 168122 734 169058 856
rect 169226 734 170162 856
rect 170330 734 171266 856
rect 171434 734 172370 856
rect 172538 734 173474 856
rect 173642 734 174578 856
rect 174746 734 175682 856
rect 175850 734 176694 856
rect 176862 734 177798 856
rect 177966 734 178902 856
rect 179070 734 180006 856
rect 180174 734 181110 856
rect 181278 734 182214 856
rect 182382 734 183318 856
rect 183486 734 184422 856
rect 184590 734 185526 856
rect 185694 734 186630 856
rect 186798 734 187734 856
rect 187902 734 188746 856
rect 188914 734 189850 856
rect 190018 734 190954 856
rect 191122 734 192058 856
rect 192226 734 193162 856
rect 193330 734 194266 856
rect 194434 734 195370 856
rect 195538 734 196474 856
rect 196642 734 197578 856
rect 197746 734 198682 856
rect 198850 734 199786 856
rect 199954 734 200798 856
rect 200966 734 201902 856
rect 202070 734 203006 856
rect 203174 734 204110 856
rect 204278 734 205214 856
rect 205382 734 206318 856
rect 206486 734 207422 856
rect 207590 734 208526 856
rect 208694 734 209630 856
rect 209798 734 210734 856
rect 210902 734 211746 856
rect 211914 734 212850 856
rect 213018 734 213954 856
rect 214122 734 215058 856
rect 215226 734 216162 856
rect 216330 734 217266 856
rect 217434 734 218370 856
rect 218538 734 219474 856
rect 219642 734 220578 856
rect 220746 734 221682 856
rect 221850 734 222786 856
rect 222954 734 223798 856
rect 223966 734 224902 856
rect 225070 734 226006 856
rect 226174 734 227110 856
rect 227278 734 228214 856
rect 228382 734 229318 856
rect 229486 734 230422 856
rect 230590 734 231526 856
rect 231694 734 232630 856
rect 232798 734 233734 856
rect 233902 734 234838 856
rect 235006 734 235850 856
rect 236018 734 236954 856
rect 237122 734 238058 856
rect 238226 734 239162 856
rect 239330 734 240266 856
rect 240434 734 241370 856
rect 241538 734 242474 856
rect 242642 734 243578 856
rect 243746 734 244682 856
rect 244850 734 245786 856
rect 245954 734 246890 856
rect 247058 734 247902 856
rect 248070 734 249006 856
rect 249174 734 250110 856
rect 250278 734 251214 856
rect 251382 734 252318 856
rect 252486 734 253422 856
rect 253590 734 254526 856
rect 254694 734 255630 856
rect 255798 734 256734 856
rect 256902 734 257838 856
rect 258006 734 258850 856
rect 259018 734 259954 856
rect 260122 734 261058 856
rect 261226 734 262162 856
rect 262330 734 263266 856
rect 263434 734 264370 856
rect 264538 734 265474 856
rect 265642 734 266578 856
rect 266746 734 267682 856
rect 267850 734 268786 856
rect 268954 734 269890 856
rect 270058 734 270902 856
rect 271070 734 272006 856
rect 272174 734 273110 856
rect 273278 734 274214 856
rect 274382 734 275318 856
rect 275486 734 276422 856
rect 276590 734 277526 856
rect 277694 734 278630 856
rect 278798 734 279734 856
rect 279902 734 280838 856
rect 281006 734 281942 856
rect 282110 734 282954 856
rect 283122 734 284058 856
rect 284226 734 285162 856
rect 285330 734 286266 856
rect 286434 734 287370 856
rect 287538 734 288474 856
rect 288642 734 289578 856
rect 289746 734 290682 856
rect 290850 734 291786 856
rect 291954 734 292890 856
rect 293058 734 293902 856
rect 294070 734 295006 856
rect 295174 734 296110 856
rect 296278 734 297214 856
rect 297382 734 298318 856
rect 298486 734 299422 856
rect 299590 734 300526 856
rect 300694 734 301630 856
rect 301798 734 302734 856
rect 302902 734 303838 856
rect 304006 734 304942 856
rect 305110 734 305954 856
rect 306122 734 307058 856
rect 307226 734 308162 856
rect 308330 734 309266 856
rect 309434 734 310370 856
rect 310538 734 311474 856
rect 311642 734 312578 856
rect 312746 734 313682 856
rect 313850 734 314786 856
rect 314954 734 315890 856
rect 316058 734 316994 856
rect 317162 734 318006 856
rect 318174 734 319110 856
rect 319278 734 320214 856
rect 320382 734 321318 856
rect 321486 734 322422 856
rect 322590 734 323526 856
rect 323694 734 324630 856
rect 324798 734 325734 856
rect 325902 734 326838 856
rect 327006 734 327942 856
rect 328110 734 329046 856
rect 329214 734 330058 856
rect 330226 734 331162 856
rect 331330 734 332266 856
rect 332434 734 333370 856
rect 333538 734 334474 856
rect 334642 734 335578 856
rect 335746 734 336682 856
rect 336850 734 337786 856
rect 337954 734 338890 856
rect 339058 734 339994 856
rect 340162 734 341006 856
rect 341174 734 342110 856
rect 342278 734 343214 856
rect 343382 734 344318 856
rect 344486 734 345422 856
rect 345590 734 346526 856
rect 346694 734 347630 856
rect 347798 734 348734 856
rect 348902 734 349838 856
rect 350006 734 350942 856
rect 351110 734 352046 856
rect 352214 734 353058 856
rect 353226 734 354162 856
rect 354330 734 355266 856
rect 355434 734 356370 856
rect 356538 734 357474 856
rect 357642 734 358578 856
rect 358746 734 359682 856
rect 359850 734 360786 856
rect 360954 734 361890 856
rect 362058 734 362994 856
rect 363162 734 364098 856
rect 364266 734 365110 856
rect 365278 734 366214 856
rect 366382 734 367318 856
rect 367486 734 368422 856
rect 368590 734 369526 856
rect 369694 734 370630 856
rect 370798 734 371734 856
rect 371902 734 372838 856
rect 373006 734 373942 856
rect 374110 734 375046 856
rect 375214 734 376058 856
rect 376226 734 377162 856
rect 377330 734 378266 856
rect 378434 734 379370 856
rect 379538 734 380474 856
rect 380642 734 381578 856
rect 381746 734 382682 856
rect 382850 734 383786 856
rect 383954 734 384890 856
rect 385058 734 385994 856
rect 386162 734 387098 856
rect 387266 734 388110 856
rect 388278 734 389214 856
rect 389382 734 390318 856
rect 390486 734 391422 856
rect 391590 734 392526 856
rect 392694 734 393630 856
rect 393798 734 394734 856
rect 394902 734 395838 856
rect 396006 734 396942 856
rect 397110 734 398046 856
rect 398214 734 399150 856
rect 399318 734 400162 856
rect 400330 734 401266 856
rect 401434 734 402370 856
rect 402538 734 403474 856
rect 403642 734 404578 856
rect 404746 734 405682 856
rect 405850 734 406786 856
rect 406954 734 407890 856
rect 408058 734 408994 856
rect 409162 734 410098 856
rect 410266 734 411202 856
rect 411370 734 412214 856
rect 412382 734 413318 856
rect 413486 734 414422 856
rect 414590 734 415526 856
rect 415694 734 416630 856
rect 416798 734 417734 856
rect 417902 734 418838 856
rect 419006 734 419942 856
rect 420110 734 421046 856
rect 421214 734 422150 856
rect 422318 734 423162 856
rect 423330 734 424266 856
rect 424434 734 425370 856
rect 425538 734 426474 856
rect 426642 734 427578 856
rect 427746 734 428682 856
rect 428850 734 429786 856
rect 429954 734 430890 856
rect 431058 734 431994 856
rect 432162 734 433098 856
rect 433266 734 434202 856
rect 434370 734 435214 856
rect 435382 734 436318 856
rect 436486 734 437422 856
rect 437590 734 438526 856
rect 438694 734 439630 856
rect 439798 734 440734 856
rect 440902 734 441838 856
rect 442006 734 442942 856
rect 443110 734 444046 856
rect 444214 734 445150 856
rect 445318 734 446254 856
rect 446422 734 447266 856
rect 447434 734 448370 856
rect 448538 734 449474 856
rect 449642 734 450578 856
rect 450746 734 451682 856
rect 451850 734 452786 856
rect 452954 734 453890 856
rect 454058 734 454994 856
rect 455162 734 456098 856
rect 456266 734 457202 856
rect 457370 734 458214 856
rect 458382 734 459318 856
rect 459486 734 460422 856
rect 460590 734 461526 856
rect 461694 734 462630 856
rect 462798 734 463734 856
rect 463902 734 464838 856
rect 465006 734 465942 856
rect 466110 734 467046 856
rect 467214 734 468150 856
rect 468318 734 469254 856
rect 469422 734 470266 856
rect 470434 734 471370 856
rect 471538 734 472474 856
rect 472642 734 473578 856
rect 473746 734 474682 856
rect 474850 734 475786 856
rect 475954 734 476890 856
rect 477058 734 477994 856
rect 478162 734 479098 856
rect 479266 734 480202 856
rect 480370 734 481306 856
rect 481474 734 482318 856
rect 482486 734 483422 856
rect 483590 734 484526 856
rect 484694 734 485630 856
rect 485798 734 486734 856
rect 486902 734 487838 856
rect 488006 734 488942 856
rect 489110 734 490046 856
rect 490214 734 491150 856
rect 491318 734 492254 856
rect 492422 734 493358 856
rect 493526 734 494370 856
rect 494538 734 495474 856
rect 495642 734 496578 856
rect 496746 734 497682 856
rect 497850 734 498786 856
rect 498954 734 499890 856
rect 500058 734 500994 856
rect 501162 734 502098 856
rect 502266 734 503202 856
rect 503370 734 504306 856
rect 504474 734 505318 856
rect 505486 734 506422 856
rect 506590 734 507526 856
rect 507694 734 508630 856
rect 508798 734 509734 856
rect 509902 734 510838 856
rect 511006 734 511942 856
rect 512110 734 513046 856
rect 513214 734 514150 856
rect 514318 734 515254 856
rect 515422 734 516358 856
rect 516526 734 517370 856
rect 517538 734 518474 856
rect 518642 734 519578 856
rect 519746 734 520682 856
rect 520850 734 521786 856
rect 521954 734 522890 856
rect 523058 734 523994 856
rect 524162 734 525098 856
rect 525266 734 526202 856
rect 526370 734 527306 856
rect 527474 734 528410 856
rect 528578 734 529422 856
rect 529590 734 530526 856
rect 530694 734 531630 856
rect 531798 734 532734 856
rect 532902 734 533838 856
rect 534006 734 534942 856
rect 535110 734 536046 856
rect 536214 734 537150 856
rect 537318 734 538254 856
rect 538422 734 539358 856
<< metal3 >>
rect 539200 309952 540000 310072
<< obsm3 >>
rect 13 2143 526768 617473
<< metal4 >>
rect 4208 2128 4528 617488
rect 19568 2128 19888 617488
rect 34928 2128 35248 617488
rect 50288 2128 50608 617488
rect 65648 2128 65968 617488
rect 81008 2128 81328 617488
rect 96368 2128 96688 617488
rect 111728 2128 112048 617488
rect 127088 2128 127408 617488
rect 142448 2128 142768 617488
rect 157808 2128 158128 617488
rect 173168 2128 173488 617488
rect 188528 2128 188848 617488
rect 203888 2128 204208 617488
rect 219248 2128 219568 617488
rect 234608 2128 234928 617488
rect 249968 2128 250288 617488
rect 265328 2128 265648 617488
rect 280688 2128 281008 617488
rect 296048 2128 296368 617488
rect 311408 2128 311728 617488
rect 326768 2128 327088 617488
rect 342128 2128 342448 617488
rect 357488 2128 357808 617488
rect 372848 2128 373168 617488
rect 388208 2128 388528 617488
rect 403568 2128 403888 617488
rect 418928 2128 419248 617488
rect 434288 2128 434608 617488
rect 449648 2128 449968 617488
rect 465008 2128 465328 617488
rect 480368 2128 480688 617488
rect 495728 2128 496048 617488
rect 511088 2128 511408 617488
rect 526448 2128 526768 617488
<< obsm4 >>
rect 19379 2347 19488 307733
rect 19968 2347 34848 307733
rect 35328 2347 50208 307733
rect 50688 2347 65568 307733
rect 66048 2347 80928 307733
rect 81408 2347 96288 307733
rect 96768 2347 111648 307733
rect 112128 2347 127008 307733
rect 127488 2347 142368 307733
rect 142848 2347 157728 307733
rect 158208 2347 173088 307733
rect 173568 2347 188448 307733
rect 188928 2347 203808 307733
rect 204288 2347 219168 307733
rect 219648 2347 234528 307733
rect 235008 2347 249888 307733
rect 250368 2347 265248 307733
rect 265728 2347 280608 307733
rect 281088 2347 284221 307733
<< labels >>
rlabel metal2 s 2318 619200 2374 620000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 143170 619200 143226 620000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 157246 619200 157302 620000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 171322 619200 171378 620000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 185398 619200 185454 620000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 199474 619200 199530 620000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 213550 619200 213606 620000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 227718 619200 227774 620000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 241794 619200 241850 620000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 255870 619200 255926 620000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 269946 619200 270002 620000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 16394 619200 16450 620000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 284022 619200 284078 620000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 298098 619200 298154 620000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 312174 619200 312230 620000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 326342 619200 326398 620000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 340418 619200 340474 620000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 354494 619200 354550 620000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 368570 619200 368626 620000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 382646 619200 382702 620000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 396722 619200 396778 620000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 410798 619200 410854 620000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 30470 619200 30526 620000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 424874 619200 424930 620000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 439042 619200 439098 620000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 453118 619200 453174 620000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 467194 619200 467250 620000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 481270 619200 481326 620000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 495346 619200 495402 620000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 509422 619200 509478 620000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 523498 619200 523554 620000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 44546 619200 44602 620000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 58622 619200 58678 620000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 72698 619200 72754 620000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 86774 619200 86830 620000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 100850 619200 100906 620000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 115018 619200 115074 620000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 129094 619200 129150 620000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 7010 619200 7066 620000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 147862 619200 147918 620000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 161938 619200 161994 620000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 176014 619200 176070 620000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 190090 619200 190146 620000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 204166 619200 204222 620000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 218334 619200 218390 620000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 232410 619200 232466 620000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 246486 619200 246542 620000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 260562 619200 260618 620000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 274638 619200 274694 620000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 21086 619200 21142 620000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 288714 619200 288770 620000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 302790 619200 302846 620000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 316866 619200 316922 620000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 331034 619200 331090 620000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 345110 619200 345166 620000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 359186 619200 359242 620000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 373262 619200 373318 620000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 387338 619200 387394 620000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 401414 619200 401470 620000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 415490 619200 415546 620000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 35162 619200 35218 620000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 429566 619200 429622 620000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 443734 619200 443790 620000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 457810 619200 457866 620000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 471886 619200 471942 620000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 485962 619200 486018 620000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 500038 619200 500094 620000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 514114 619200 514170 620000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 528190 619200 528246 620000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 49238 619200 49294 620000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 63314 619200 63370 620000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 77390 619200 77446 620000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 91466 619200 91522 620000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 105542 619200 105598 620000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 119710 619200 119766 620000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 133786 619200 133842 620000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 11702 619200 11758 620000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 152554 619200 152610 620000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 166630 619200 166686 620000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 180706 619200 180762 620000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 194782 619200 194838 620000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 208858 619200 208914 620000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 223026 619200 223082 620000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 237102 619200 237158 620000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 251178 619200 251234 620000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 265254 619200 265310 620000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 279330 619200 279386 620000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 25778 619200 25834 620000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 293406 619200 293462 620000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 307482 619200 307538 620000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 321558 619200 321614 620000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 335726 619200 335782 620000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 349802 619200 349858 620000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 363878 619200 363934 620000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 377954 619200 378010 620000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 392030 619200 392086 620000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 406106 619200 406162 620000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 420182 619200 420238 620000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 39854 619200 39910 620000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 434350 619200 434406 620000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 448426 619200 448482 620000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 462502 619200 462558 620000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 476578 619200 476634 620000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 490654 619200 490710 620000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 504730 619200 504786 620000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 518806 619200 518862 620000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 532882 619200 532938 620000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 53930 619200 53986 620000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 68006 619200 68062 620000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 82082 619200 82138 620000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 96158 619200 96214 620000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 110326 619200 110382 620000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 124402 619200 124458 620000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 138478 619200 138534 620000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 537206 0 537262 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 538310 0 538366 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 539414 0 539470 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 445206 0 445262 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 448426 0 448482 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 451738 0 451794 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 455050 0 455106 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 458270 0 458326 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 461582 0 461638 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 464894 0 464950 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 468206 0 468262 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 471426 0 471482 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 474738 0 474794 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 478050 0 478106 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 481362 0 481418 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 484582 0 484638 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 487894 0 487950 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 491206 0 491262 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 494426 0 494482 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 497738 0 497794 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 501050 0 501106 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 504362 0 504418 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 507582 0 507638 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 510894 0 510950 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 514206 0 514262 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 517426 0 517482 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 520738 0 520794 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 524050 0 524106 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 527362 0 527418 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 530582 0 530638 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 533894 0 533950 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 218426 0 218482 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 238114 0 238170 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 241426 0 241482 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 247958 0 248014 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 251270 0 251326 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 254582 0 254638 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 264426 0 264482 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 270958 0 271014 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 280894 0 280950 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 284114 0 284170 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 290738 0 290794 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 297270 0 297326 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 303894 0 303950 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 307114 0 307170 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 313738 0 313794 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 317050 0 317106 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 320270 0 320326 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 323582 0 323638 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 326894 0 326950 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 333426 0 333482 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 336738 0 336794 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 343270 0 343326 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 349894 0 349950 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 353114 0 353170 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 356426 0 356482 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 359738 0 359794 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 363050 0 363106 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 366270 0 366326 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 369582 0 369638 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 372894 0 372950 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 376114 0 376170 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 379426 0 379482 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 382738 0 382794 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 386050 0 386106 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 389270 0 389326 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 392582 0 392638 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 395894 0 395950 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 399206 0 399262 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 402426 0 402482 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 405738 0 405794 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 409050 0 409106 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 412270 0 412326 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 415582 0 415638 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 418894 0 418950 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 422206 0 422262 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 425426 0 425482 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 428738 0 428794 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 432050 0 432106 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 435270 0 435326 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 438582 0 438638 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 441894 0 441950 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 446310 0 446366 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 449530 0 449586 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 452842 0 452898 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 456154 0 456210 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 459374 0 459430 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 462686 0 462742 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 465998 0 466054 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 469310 0 469366 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 472530 0 472586 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 475842 0 475898 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 479154 0 479210 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 482374 0 482430 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 485686 0 485742 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 488998 0 489054 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 492310 0 492366 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 495530 0 495586 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 498842 0 498898 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 502154 0 502210 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 505374 0 505430 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 508686 0 508742 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 511998 0 512054 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 515310 0 515366 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 518530 0 518586 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 521842 0 521898 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 525154 0 525210 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 528466 0 528522 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 531686 0 531742 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 534998 0 535054 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 170218 0 170274 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 180062 0 180118 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 196530 0 196586 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 199842 0 199898 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 203062 0 203118 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 206374 0 206430 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 209686 0 209742 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 216218 0 216274 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 219530 0 219586 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 229374 0 229430 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 232686 0 232742 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 235906 0 235962 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 242530 0 242586 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 245842 0 245898 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 252374 0 252430 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 255686 0 255742 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 262218 0 262274 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 265530 0 265586 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 272062 0 272118 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 275374 0 275430 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 281998 0 282054 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 285218 0 285274 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 288530 0 288586 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 291842 0 291898 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 295062 0 295118 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 298374 0 298430 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 301686 0 301742 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 304998 0 305054 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 308218 0 308274 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 311530 0 311586 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 314842 0 314898 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 318062 0 318118 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 321374 0 321430 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 324686 0 324742 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 327998 0 328054 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 331218 0 331274 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 334530 0 334586 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 337842 0 337898 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 341062 0 341118 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 344374 0 344430 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 137374 0 137430 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 347686 0 347742 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 350998 0 351054 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 354218 0 354274 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 357530 0 357586 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 360842 0 360898 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 364154 0 364210 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 367374 0 367430 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 370686 0 370742 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 373998 0 374054 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 377218 0 377274 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 380530 0 380586 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 383842 0 383898 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 387154 0 387210 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 390374 0 390430 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 393686 0 393742 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 396998 0 397054 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 400218 0 400274 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 403530 0 403586 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 406842 0 406898 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 410154 0 410210 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 413374 0 413430 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 416686 0 416742 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 419998 0 420054 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 423218 0 423274 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 426530 0 426586 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 429842 0 429898 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 433154 0 433210 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 436374 0 436430 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 439686 0 439742 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 442998 0 443054 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 447322 0 447378 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 450634 0 450690 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 453946 0 454002 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 457258 0 457314 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 460478 0 460534 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 463790 0 463846 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 467102 0 467158 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 470322 0 470378 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 473634 0 473690 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 476946 0 477002 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 480258 0 480314 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 483478 0 483534 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 486790 0 486846 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 490102 0 490158 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 493414 0 493470 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 496634 0 496690 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 499946 0 500002 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 503258 0 503314 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 506478 0 506534 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 509790 0 509846 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 513102 0 513158 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 516414 0 516470 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 519634 0 519690 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 522946 0 523002 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 526258 0 526314 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 529478 0 529534 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 532790 0 532846 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 536102 0 536158 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 204166 0 204222 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 230478 0 230534 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 240322 0 240378 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 246946 0 247002 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 260010 0 260066 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 263322 0 263378 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 266634 0 266690 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 269946 0 270002 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 273166 0 273222 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 276478 0 276534 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 279790 0 279846 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 286322 0 286378 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 289634 0 289690 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 292946 0 293002 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 296166 0 296222 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 306010 0 306066 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 309322 0 309378 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 312634 0 312690 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 315946 0 316002 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 319166 0 319222 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 322478 0 322534 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 325790 0 325846 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 329102 0 329158 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 335634 0 335690 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 338946 0 339002 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 342166 0 342222 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 345478 0 345534 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 348790 0 348846 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 352102 0 352158 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 355322 0 355378 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 358634 0 358690 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 361946 0 362002 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 365166 0 365222 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 368478 0 368534 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 371790 0 371846 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 375102 0 375158 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 378322 0 378378 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 381634 0 381690 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 384946 0 385002 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 388166 0 388222 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 391478 0 391534 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 394790 0 394846 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 398102 0 398158 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 401322 0 401378 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 404634 0 404690 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 407946 0 408002 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 411258 0 411314 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 414478 0 414534 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 417790 0 417846 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 421102 0 421158 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 424322 0 424378 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 430946 0 431002 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 434258 0 434314 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 437478 0 437534 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 440790 0 440846 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 444102 0 444158 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 617488 6 vccd1
port 502 nsew power bidirectional
rlabel metal2 s 537574 619200 537630 620000 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 617488 6 vssd1
port 504 nsew ground bidirectional
rlabel metal3 s 539200 309952 540000 310072 6 vssd1
port 505 nsew ground bidirectional
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 506 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 507 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_ack_o
port 508 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[0]
port 509 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_adr_i[10]
port 510 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_adr_i[11]
port 511 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_adr_i[12]
port 512 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_adr_i[13]
port 513 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_adr_i[14]
port 514 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_adr_i[15]
port 515 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 wbs_adr_i[16]
port 516 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wbs_adr_i[17]
port 517 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wbs_adr_i[18]
port 518 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[19]
port 519 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[1]
port 520 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 wbs_adr_i[20]
port 521 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 wbs_adr_i[21]
port 522 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 wbs_adr_i[22]
port 523 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_adr_i[23]
port 524 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 wbs_adr_i[24]
port 525 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 wbs_adr_i[25]
port 526 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 wbs_adr_i[26]
port 527 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 wbs_adr_i[27]
port 528 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 wbs_adr_i[28]
port 529 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 wbs_adr_i[29]
port 530 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[2]
port 531 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 wbs_adr_i[30]
port 532 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 wbs_adr_i[31]
port 533 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[3]
port 534 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[4]
port 535 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[5]
port 536 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[6]
port 537 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[7]
port 538 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[8]
port 539 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_adr_i[9]
port 540 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_cyc_i
port 541 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[0]
port 542 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[10]
port 543 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_i[11]
port 544 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_i[12]
port 545 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_i[13]
port 546 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_i[14]
port 547 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[15]
port 548 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_dat_i[16]
port 549 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_i[17]
port 550 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_i[18]
port 551 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 wbs_dat_i[19]
port 552 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[1]
port 553 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_i[20]
port 554 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_i[21]
port 555 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[22]
port 556 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 wbs_dat_i[23]
port 557 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 wbs_dat_i[24]
port 558 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 wbs_dat_i[25]
port 559 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 wbs_dat_i[26]
port 560 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 wbs_dat_i[27]
port 561 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 wbs_dat_i[28]
port 562 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 wbs_dat_i[29]
port 563 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[2]
port 564 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 wbs_dat_i[30]
port 565 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 wbs_dat_i[31]
port 566 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[3]
port 567 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[4]
port 568 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[5]
port 569 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[6]
port 570 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[7]
port 571 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[8]
port 572 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_i[9]
port 573 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[0]
port 574 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_o[10]
port 575 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[11]
port 576 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[12]
port 577 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[13]
port 578 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_o[14]
port 579 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_o[15]
port 580 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_o[16]
port 581 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 wbs_dat_o[17]
port 582 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_o[18]
port 583 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 wbs_dat_o[19]
port 584 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[1]
port 585 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 wbs_dat_o[20]
port 586 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 wbs_dat_o[21]
port 587 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 wbs_dat_o[22]
port 588 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[23]
port 589 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[24]
port 590 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[25]
port 591 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_o[26]
port 592 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 wbs_dat_o[27]
port 593 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_o[28]
port 594 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 wbs_dat_o[29]
port 595 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[2]
port 596 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 wbs_dat_o[30]
port 597 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 wbs_dat_o[31]
port 598 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_o[3]
port 599 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[4]
port 600 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_o[5]
port 601 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[6]
port 602 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[7]
port 603 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[8]
port 604 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 wbs_dat_o[9]
port 605 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_sel_i[0]
port 606 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_sel_i[1]
port 607 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_sel_i[2]
port 608 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_sel_i[3]
port 609 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_stb_i
port 610 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_we_i
port 611 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 540000 620000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 215875434
string GDS_FILE /home/asic/mont/SonarOnChip8/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 1646940
<< end >>

